module rotate_lut (
    input logic [9:0] counter,        // Counter ranging from 0 to 783
    output logic [9:0] rot_addr       // Rotated address output
);

    always_comb begin
	  case (counter) 
	    10'b0: rot_addr = 10'b0;
	    10'b1: rot_addr = 10'b0;
	    10'b10: rot_addr = 10'b0;
	    10'b11: rot_addr = 10'b0;
	    10'b100: rot_addr = 10'b0;
	    10'b101: rot_addr = 10'b0;
	    10'b110: rot_addr = 10'b0;
	    10'b111: rot_addr = 10'b0;
	    10'b1000: rot_addr = 10'b0;
	    10'b1001: rot_addr = 10'b0;
	    10'b1010: rot_addr = 10'b0;
	    10'b1011: rot_addr = 10'b10000;
	    10'b1100: rot_addr = 10'b10001;
	    10'b1101: rot_addr = 10'b101110;
	    10'b1110: rot_addr = 10'b101111;
	    10'b1111: rot_addr = 10'b110000;
	    10'b10000: rot_addr = 10'b1001101;
	    10'b10001: rot_addr = 10'b1001110;
	    10'b10010: rot_addr = 10'b1001111;
	    10'b10011: rot_addr = 10'b1101011;
	    10'b10100: rot_addr = 10'b1101100;
	    10'b10101: rot_addr = 10'b1101101;
	    10'b10110: rot_addr = 10'b10001010;
	    10'b10111: rot_addr = 10'b10001011;
	    10'b11000: rot_addr = 10'b10001100;
	    10'b11001: rot_addr = 10'b0;
	    10'b11010: rot_addr = 10'b0;
	    10'b11011: rot_addr = 10'b0;
	    10'b11100: rot_addr = 10'b0;
	    10'b11101: rot_addr = 10'b0;
	    10'b11110: rot_addr = 10'b0;
	    10'b11111: rot_addr = 10'b0;
	    10'b100000: rot_addr = 10'b0;
	    10'b100001: rot_addr = 10'b0;
	    10'b100010: rot_addr = 10'b0;
	    10'b100011: rot_addr = 10'b0;
	    10'b100100: rot_addr = 10'b1101;
	    10'b100101: rot_addr = 10'b1110;
	    10'b100110: rot_addr = 10'b1111;
	    10'b100111: rot_addr = 10'b101100;
	    10'b101000: rot_addr = 10'b101101;
	    10'b101001: rot_addr = 10'b101110;
	    10'b101010: rot_addr = 10'b1001010;
	    10'b101011: rot_addr = 10'b1001011;
	    10'b101100: rot_addr = 10'b1001100;
	    10'b101101: rot_addr = 10'b1101001;
	    10'b101110: rot_addr = 10'b1101010;
	    10'b101111: rot_addr = 10'b1101011;
	    10'b110000: rot_addr = 10'b10001000;
	    10'b110001: rot_addr = 10'b10001001;
	    10'b110010: rot_addr = 10'b10100110;
	    10'b110011: rot_addr = 10'b10100111;
	    10'b110100: rot_addr = 10'b10101000;
	    10'b110101: rot_addr = 10'b0;
	    10'b110110: rot_addr = 10'b0;
	    10'b110111: rot_addr = 10'b0;
	    10'b111000: rot_addr = 10'b0;
	    10'b111001: rot_addr = 10'b0;
	    10'b111010: rot_addr = 10'b0;
	    10'b111011: rot_addr = 10'b0;
	    10'b111100: rot_addr = 10'b0;
	    10'b111101: rot_addr = 10'b1010;
	    10'b111110: rot_addr = 10'b1011;
	    10'b111111: rot_addr = 10'b1100;
	    10'b1000000: rot_addr = 10'b101000;
	    10'b1000001: rot_addr = 10'b101001;
	    10'b1000010: rot_addr = 10'b101010;
	    10'b1000011: rot_addr = 10'b1000111;
	    10'b1000100: rot_addr = 10'b1001000;
	    10'b1000101: rot_addr = 10'b1001001;
	    10'b1000110: rot_addr = 10'b1100110;
	    10'b1000111: rot_addr = 10'b1100111;
	    10'b1001000: rot_addr = 10'b1101000;
	    10'b1001001: rot_addr = 10'b10000101;
	    10'b1001010: rot_addr = 10'b10000110;
	    10'b1001011: rot_addr = 10'b10000111;
	    10'b1001100: rot_addr = 10'b10100100;
	    10'b1001101: rot_addr = 10'b10100101;
	    10'b1001110: rot_addr = 10'b10100110;
	    10'b1001111: rot_addr = 10'b11000011;
	    10'b1010000: rot_addr = 10'b11000100;
	    10'b1010001: rot_addr = 10'b11000100;
	    10'b1010010: rot_addr = 10'b0;
	    10'b1010011: rot_addr = 10'b0;
	    10'b1010100: rot_addr = 10'b0;
	    10'b1010101: rot_addr = 10'b0;
	    10'b1010110: rot_addr = 10'b110;
	    10'b1010111: rot_addr = 10'b111;
	    10'b1011000: rot_addr = 10'b1000;
	    10'b1011001: rot_addr = 10'b100101;
	    10'b1011010: rot_addr = 10'b100110;
	    10'b1011011: rot_addr = 10'b100111;
	    10'b1011100: rot_addr = 10'b1000100;
	    10'b1011101: rot_addr = 10'b1000101;
	    10'b1011110: rot_addr = 10'b1000110;
	    10'b1011111: rot_addr = 10'b1100011;
	    10'b1100000: rot_addr = 10'b1100100;
	    10'b1100001: rot_addr = 10'b1100101;
	    10'b1100010: rot_addr = 10'b10000010;
	    10'b1100011: rot_addr = 10'b10000011;
	    10'b1100100: rot_addr = 10'b10000100;
	    10'b1100101: rot_addr = 10'b10100001;
	    10'b1100110: rot_addr = 10'b10100010;
	    10'b1100111: rot_addr = 10'b10100010;
	    10'b1101000: rot_addr = 10'b10111111;
	    10'b1101001: rot_addr = 10'b11000000;
	    10'b1101010: rot_addr = 10'b11000001;
	    10'b1101011: rot_addr = 10'b11011110;
	    10'b1101100: rot_addr = 10'b11011111;
	    10'b1101101: rot_addr = 10'b11100000;
	    10'b1101110: rot_addr = 10'b0;
	    10'b1101111: rot_addr = 10'b0;
	    10'b1110000: rot_addr = 10'b100;
	    10'b1110001: rot_addr = 10'b101;
	    10'b1110010: rot_addr = 10'b110;
	    10'b1110011: rot_addr = 10'b100011;
	    10'b1110100: rot_addr = 10'b100100;
	    10'b1110101: rot_addr = 10'b1000001;
	    10'b1110110: rot_addr = 10'b1000010;
	    10'b1110111: rot_addr = 10'b1000011;
	    10'b1111000: rot_addr = 10'b1100000;
	    10'b1111001: rot_addr = 10'b1100001;
	    10'b1111010: rot_addr = 10'b1100010;
	    10'b1111011: rot_addr = 10'b1111111;
	    10'b1111100: rot_addr = 10'b10000000;
	    10'b1111101: rot_addr = 10'b10000000;
	    10'b1111110: rot_addr = 10'b10011101;
	    10'b1111111: rot_addr = 10'b10011110;
	    10'b10000000: rot_addr = 10'b10011111;
	    10'b10000001: rot_addr = 10'b10111100;
	    10'b10000010: rot_addr = 10'b10111101;
	    10'b10000011: rot_addr = 10'b10111110;
	    10'b10000100: rot_addr = 10'b11011011;
	    10'b10000101: rot_addr = 10'b11011100;
	    10'b10000110: rot_addr = 10'b11011101;
	    10'b10000111: rot_addr = 10'b11111010;
	    10'b10001000: rot_addr = 10'b11111011;
	    10'b10001001: rot_addr = 10'b11111100;
	    10'b10001010: rot_addr = 10'b0;
	    10'b10001011: rot_addr = 10'b0;
	    10'b10001100: rot_addr = 10'b100000;
	    10'b10001101: rot_addr = 10'b100001;
	    10'b10001110: rot_addr = 10'b100010;
	    10'b10001111: rot_addr = 10'b111111;
	    10'b10010000: rot_addr = 10'b1000000;
	    10'b10010001: rot_addr = 10'b1000001;
	    10'b10010010: rot_addr = 10'b1011110;
	    10'b10010011: rot_addr = 10'b1011111;
	    10'b10010100: rot_addr = 10'b1011111;
	    10'b10010101: rot_addr = 10'b1111100;
	    10'b10010110: rot_addr = 10'b1111101;
	    10'b10010111: rot_addr = 10'b10011010;
	    10'b10011000: rot_addr = 10'b10011011;
	    10'b10011001: rot_addr = 10'b10011100;
	    10'b10011010: rot_addr = 10'b10111001;
	    10'b10011011: rot_addr = 10'b10111010;
	    10'b10011100: rot_addr = 10'b10111011;
	    10'b10011101: rot_addr = 10'b11011000;
	    10'b10011110: rot_addr = 10'b11011001;
	    10'b10011111: rot_addr = 10'b11011010;
	    10'b10100000: rot_addr = 10'b11110111;
	    10'b10100001: rot_addr = 10'b11111000;
	    10'b10100010: rot_addr = 10'b11111001;
	    10'b10100011: rot_addr = 10'b100010110;
	    10'b10100100: rot_addr = 10'b100010110;
	    10'b10100101: rot_addr = 10'b100010111;
	    10'b10100110: rot_addr = 10'b100110100;
	    10'b10100111: rot_addr = 10'b0;
	    10'b10101000: rot_addr = 10'b111100;
	    10'b10101001: rot_addr = 10'b111101;
	    10'b10101010: rot_addr = 10'b111101;
	    10'b10101011: rot_addr = 10'b1011010;
	    10'b10101100: rot_addr = 10'b1011011;
	    10'b10101101: rot_addr = 10'b1011100;
	    10'b10101110: rot_addr = 10'b1111001;
	    10'b10101111: rot_addr = 10'b1111010;
	    10'b10110000: rot_addr = 10'b1111011;
	    10'b10110001: rot_addr = 10'b10011000;
	    10'b10110010: rot_addr = 10'b10011001;
	    10'b10110011: rot_addr = 10'b10011010;
	    10'b10110100: rot_addr = 10'b10110111;
	    10'b10110101: rot_addr = 10'b10111000;
	    10'b10110110: rot_addr = 10'b10111001;
	    10'b10110111: rot_addr = 10'b11010110;
	    10'b10111000: rot_addr = 10'b11010111;
	    10'b10111001: rot_addr = 10'b11110100;
	    10'b10111010: rot_addr = 10'b11110100;
	    10'b10111011: rot_addr = 10'b11110101;
	    10'b10111100: rot_addr = 10'b100010010;
	    10'b10111101: rot_addr = 10'b100010011;
	    10'b10111110: rot_addr = 10'b100010100;
	    10'b10111111: rot_addr = 10'b100110001;
	    10'b11000000: rot_addr = 10'b100110010;
	    10'b11000001: rot_addr = 10'b100110011;
	    10'b11000010: rot_addr = 10'b101010000;
	    10'b11000011: rot_addr = 10'b0;
	    10'b11000100: rot_addr = 10'b1010111;
	    10'b11000101: rot_addr = 10'b1011000;
	    10'b11000110: rot_addr = 10'b1011001;
	    10'b11000111: rot_addr = 10'b1110110;
	    10'b11001000: rot_addr = 10'b1110111;
	    10'b11001001: rot_addr = 10'b1111000;
	    10'b11001010: rot_addr = 10'b10010101;
	    10'b11001011: rot_addr = 10'b10010110;
	    10'b11001100: rot_addr = 10'b10010111;
	    10'b11001101: rot_addr = 10'b10110100;
	    10'b11001110: rot_addr = 10'b10110101;
	    10'b11001111: rot_addr = 10'b10110110;
	    10'b11010000: rot_addr = 10'b11010011;
	    10'b11010001: rot_addr = 10'b11010011;
	    10'b11010010: rot_addr = 10'b11010100;
	    10'b11010011: rot_addr = 10'b11110001;
	    10'b11010100: rot_addr = 10'b11110010;
	    10'b11010101: rot_addr = 10'b11110011;
	    10'b11010110: rot_addr = 10'b100010000;
	    10'b11010111: rot_addr = 10'b100010001;
	    10'b11011000: rot_addr = 10'b100010010;
	    10'b11011001: rot_addr = 10'b100101111;
	    10'b11011010: rot_addr = 10'b100110000;
	    10'b11011011: rot_addr = 10'b101001101;
	    10'b11011100: rot_addr = 10'b101001110;
	    10'b11011101: rot_addr = 10'b101001111;
	    10'b11011110: rot_addr = 10'b101101100;
	    10'b11011111: rot_addr = 10'b0;
	    10'b11100000: rot_addr = 10'b1110011;
	    10'b11100001: rot_addr = 10'b1110100;
	    10'b11100010: rot_addr = 10'b1110101;
	    10'b11100011: rot_addr = 10'b10010010;
	    10'b11100100: rot_addr = 10'b10010011;
	    10'b11100101: rot_addr = 10'b10010100;
	    10'b11100110: rot_addr = 10'b10110001;
	    10'b11100111: rot_addr = 10'b10110001;
	    10'b11101000: rot_addr = 10'b10110010;
	    10'b11101001: rot_addr = 10'b11001111;
	    10'b11101010: rot_addr = 10'b11010000;
	    10'b11101011: rot_addr = 10'b11010001;
	    10'b11101100: rot_addr = 10'b11101110;
	    10'b11101101: rot_addr = 10'b11101111;
	    10'b11101110: rot_addr = 10'b11110000;
	    10'b11101111: rot_addr = 10'b100001101;
	    10'b11110000: rot_addr = 10'b100001110;
	    10'b11110001: rot_addr = 10'b100001111;
	    10'b11110010: rot_addr = 10'b100101100;
	    10'b11110011: rot_addr = 10'b100101101;
	    10'b11110100: rot_addr = 10'b100101110;
	    10'b11110101: rot_addr = 10'b101001011;
	    10'b11110110: rot_addr = 10'b101001100;
	    10'b11110111: rot_addr = 10'b101001101;
	    10'b11111000: rot_addr = 10'b101101001;
	    10'b11111001: rot_addr = 10'b101101010;
	    10'b11111010: rot_addr = 10'b101101011;
	    10'b11111011: rot_addr = 10'b110001000;
	    10'b11111100: rot_addr = 10'b10001111;
	    10'b11111101: rot_addr = 10'b10001111;
	    10'b11111110: rot_addr = 10'b10010000;
	    10'b11111111: rot_addr = 10'b10101101;
	    10'b100000000: rot_addr = 10'b10101110;
	    10'b100000001: rot_addr = 10'b10101111;
	    10'b100000010: rot_addr = 10'b11001100;
	    10'b100000011: rot_addr = 10'b11001101;
	    10'b100000100: rot_addr = 10'b11001110;
	    10'b100000101: rot_addr = 10'b11101011;
	    10'b100000110: rot_addr = 10'b11101100;
	    10'b100000111: rot_addr = 10'b11101101;
	    10'b100001000: rot_addr = 10'b100001010;
	    10'b100001001: rot_addr = 10'b100001011;
	    10'b100001010: rot_addr = 10'b100001100;
	    10'b100001011: rot_addr = 10'b100101001;
	    10'b100001100: rot_addr = 10'b100101010;
	    10'b100001101: rot_addr = 10'b100101011;
	    10'b100001110: rot_addr = 10'b101000111;
	    10'b100001111: rot_addr = 10'b101001000;
	    10'b100010000: rot_addr = 10'b101001001;
	    10'b100010001: rot_addr = 10'b101100110;
	    10'b100010010: rot_addr = 10'b101100111;
	    10'b100010011: rot_addr = 10'b101101000;
	    10'b100010100: rot_addr = 10'b110000101;
	    10'b100010101: rot_addr = 10'b110000110;
	    10'b100010110: rot_addr = 10'b110000111;
	    10'b100010111: rot_addr = 10'b110100100;
	    10'b100011000: rot_addr = 10'b10001110;
	    10'b100011001: rot_addr = 10'b10101011;
	    10'b100011010: rot_addr = 10'b10101100;
	    10'b100011011: rot_addr = 10'b10101101;
	    10'b100011100: rot_addr = 10'b11001010;
	    10'b100011101: rot_addr = 10'b11001011;
	    10'b100011110: rot_addr = 10'b11101000;
	    10'b100011111: rot_addr = 10'b11101001;
	    10'b100100000: rot_addr = 10'b11101010;
	    10'b100100001: rot_addr = 10'b100000111;
	    10'b100100010: rot_addr = 10'b100001000;
	    10'b100100011: rot_addr = 10'b100001001;
	    10'b100100100: rot_addr = 10'b100100101;
	    10'b100100101: rot_addr = 10'b100100110;
	    10'b100100110: rot_addr = 10'b100100111;
	    10'b100100111: rot_addr = 10'b101000100;
	    10'b100101000: rot_addr = 10'b101000101;
	    10'b100101001: rot_addr = 10'b101000110;
	    10'b100101010: rot_addr = 10'b101100011;
	    10'b100101011: rot_addr = 10'b101100100;
	    10'b100101100: rot_addr = 10'b101100101;
	    10'b100101101: rot_addr = 10'b110000010;
	    10'b100101110: rot_addr = 10'b110000011;
	    10'b100101111: rot_addr = 10'b110000100;
	    10'b100110000: rot_addr = 10'b110100001;
	    10'b100110001: rot_addr = 10'b110100010;
	    10'b100110010: rot_addr = 10'b110100011;
	    10'b100110011: rot_addr = 10'b111000000;
	    10'b100110100: rot_addr = 10'b10101010;
	    10'b100110101: rot_addr = 10'b11000111;
	    10'b100110110: rot_addr = 10'b11001000;
	    10'b100110111: rot_addr = 10'b11001001;
	    10'b100111000: rot_addr = 10'b11100110;
	    10'b100111001: rot_addr = 10'b11100111;
	    10'b100111010: rot_addr = 10'b11101000;
	    10'b100111011: rot_addr = 10'b100000100;
	    10'b100111100: rot_addr = 10'b100000101;
	    10'b100111101: rot_addr = 10'b100000110;
	    10'b100111110: rot_addr = 10'b100100011;
	    10'b100111111: rot_addr = 10'b100100100;
	    10'b101000000: rot_addr = 10'b100100101;
	    10'b101000001: rot_addr = 10'b101000010;
	    10'b101000010: rot_addr = 10'b101000011;
	    10'b101000011: rot_addr = 10'b101100000;
	    10'b101000100: rot_addr = 10'b101100001;
	    10'b101000101: rot_addr = 10'b101100010;
	    10'b101000110: rot_addr = 10'b101111111;
	    10'b101000111: rot_addr = 10'b110000000;
	    10'b101001000: rot_addr = 10'b110000001;
	    10'b101001001: rot_addr = 10'b110011110;
	    10'b101001010: rot_addr = 10'b110011111;
	    10'b101001011: rot_addr = 10'b110011111;
	    10'b101001100: rot_addr = 10'b110111100;
	    10'b101001101: rot_addr = 10'b110111101;
	    10'b101001110: rot_addr = 10'b110111110;
	    10'b101001111: rot_addr = 10'b111011011;
	    10'b101010000: rot_addr = 10'b11000110;
	    10'b101010001: rot_addr = 10'b11100010;
	    10'b101010010: rot_addr = 10'b11100011;
	    10'b101010011: rot_addr = 10'b11100100;
	    10'b101010100: rot_addr = 10'b100000001;
	    10'b101010101: rot_addr = 10'b100000010;
	    10'b101010110: rot_addr = 10'b100000011;
	    10'b101010111: rot_addr = 10'b100100000;
	    10'b101011000: rot_addr = 10'b100100001;
	    10'b101011001: rot_addr = 10'b100100010;
	    10'b101011010: rot_addr = 10'b100111111;
	    10'b101011011: rot_addr = 10'b101000000;
	    10'b101011100: rot_addr = 10'b101000001;
	    10'b101011101: rot_addr = 10'b101011110;
	    10'b101011110: rot_addr = 10'b101011111;
	    10'b101011111: rot_addr = 10'b101100000;
	    10'b101100000: rot_addr = 10'b101111101;
	    10'b101100001: rot_addr = 10'b101111110;
	    10'b101100010: rot_addr = 10'b101111110;
	    10'b101100011: rot_addr = 10'b110011011;
	    10'b101100100: rot_addr = 10'b110011100;
	    10'b101100101: rot_addr = 10'b110111001;
	    10'b101100110: rot_addr = 10'b110111010;
	    10'b101100111: rot_addr = 10'b110111011;
	    10'b101101000: rot_addr = 10'b111011000;
	    10'b101101001: rot_addr = 10'b111011001;
	    10'b101101010: rot_addr = 10'b111011010;
	    10'b101101011: rot_addr = 10'b111110111;
	    10'b101101100: rot_addr = 10'b11100001;
	    10'b101101101: rot_addr = 10'b11111110;
	    10'b101101110: rot_addr = 10'b11111111;
	    10'b101101111: rot_addr = 10'b100000000;
	    10'b101110000: rot_addr = 10'b100011101;
	    10'b101110001: rot_addr = 10'b100011110;
	    10'b101110010: rot_addr = 10'b100011111;
	    10'b101110011: rot_addr = 10'b100111100;
	    10'b101110100: rot_addr = 10'b100111101;
	    10'b101110101: rot_addr = 10'b100111110;
	    10'b101110110: rot_addr = 10'b101011011;
	    10'b101110111: rot_addr = 10'b101011100;
	    10'b101111000: rot_addr = 10'b101011100;
	    10'b101111001: rot_addr = 10'b101111001;
	    10'b101111010: rot_addr = 10'b101111010;
	    10'b101111011: rot_addr = 10'b101111011;
	    10'b101111100: rot_addr = 10'b110011000;
	    10'b101111101: rot_addr = 10'b110011001;
	    10'b101111110: rot_addr = 10'b110011010;
	    10'b101111111: rot_addr = 10'b110110111;
	    10'b110000000: rot_addr = 10'b110111000;
	    10'b110000001: rot_addr = 10'b110111001;
	    10'b110000010: rot_addr = 10'b111010110;
	    10'b110000011: rot_addr = 10'b111010111;
	    10'b110000100: rot_addr = 10'b111011000;
	    10'b110000101: rot_addr = 10'b111110101;
	    10'b110000110: rot_addr = 10'b111110110;
	    10'b110000111: rot_addr = 10'b1000010011;
	    10'b110001000: rot_addr = 10'b11111101;
	    10'b110001001: rot_addr = 10'b100011010;
	    10'b110001010: rot_addr = 10'b100011011;
	    10'b110001011: rot_addr = 10'b100011100;
	    10'b110001100: rot_addr = 10'b100111001;
	    10'b110001101: rot_addr = 10'b100111010;
	    10'b110001110: rot_addr = 10'b100111010;
	    10'b110001111: rot_addr = 10'b101010111;
	    10'b110010000: rot_addr = 10'b101011000;
	    10'b110010001: rot_addr = 10'b101011001;
	    10'b110010010: rot_addr = 10'b101110110;
	    10'b110010011: rot_addr = 10'b101110111;
	    10'b110010100: rot_addr = 10'b101111000;
	    10'b110010101: rot_addr = 10'b110010101;
	    10'b110010110: rot_addr = 10'b110010110;
	    10'b110010111: rot_addr = 10'b110010111;
	    10'b110011000: rot_addr = 10'b110110100;
	    10'b110011001: rot_addr = 10'b110110101;
	    10'b110011010: rot_addr = 10'b110110110;
	    10'b110011011: rot_addr = 10'b111010011;
	    10'b110011100: rot_addr = 10'b111010100;
	    10'b110011101: rot_addr = 10'b111010101;
	    10'b110011110: rot_addr = 10'b111110010;
	    10'b110011111: rot_addr = 10'b111110010;
	    10'b110100000: rot_addr = 10'b111110011;
	    10'b110100001: rot_addr = 10'b1000010000;
	    10'b110100010: rot_addr = 10'b1000010001;
	    10'b110100011: rot_addr = 10'b1000010010;
	    10'b110100100: rot_addr = 10'b100011001;
	    10'b110100101: rot_addr = 10'b100011001;
	    10'b110100110: rot_addr = 10'b100110110;
	    10'b110100111: rot_addr = 10'b100110111;
	    10'b110101000: rot_addr = 10'b101010100;
	    10'b110101001: rot_addr = 10'b101010101;
	    10'b110101010: rot_addr = 10'b101010110;
	    10'b110101011: rot_addr = 10'b101110011;
	    10'b110101100: rot_addr = 10'b101110100;
	    10'b110101101: rot_addr = 10'b101110101;
	    10'b110101110: rot_addr = 10'b110010010;
	    10'b110101111: rot_addr = 10'b110010011;
	    10'b110110000: rot_addr = 10'b110010100;
	    10'b110110001: rot_addr = 10'b110110001;
	    10'b110110010: rot_addr = 10'b110110010;
	    10'b110110011: rot_addr = 10'b110110011;
	    10'b110110100: rot_addr = 10'b111010000;
	    10'b110110101: rot_addr = 10'b111010000;
	    10'b110110110: rot_addr = 10'b111010001;
	    10'b110110111: rot_addr = 10'b111101110;
	    10'b110111000: rot_addr = 10'b111101111;
	    10'b110111001: rot_addr = 10'b111110000;
	    10'b110111010: rot_addr = 10'b1000001101;
	    10'b110111011: rot_addr = 10'b1000001110;
	    10'b110111100: rot_addr = 10'b1000001111;
	    10'b110111101: rot_addr = 10'b1000101100;
	    10'b110111110: rot_addr = 10'b1000101101;
	    10'b110111111: rot_addr = 10'b1000101110;
	    10'b111000000: rot_addr = 10'b0;
	    10'b111000001: rot_addr = 10'b100110101;
	    10'b111000010: rot_addr = 10'b101010010;
	    10'b111000011: rot_addr = 10'b101010011;
	    10'b111000100: rot_addr = 10'b101010100;
	    10'b111000101: rot_addr = 10'b101110001;
	    10'b111000110: rot_addr = 10'b101110010;
	    10'b111000111: rot_addr = 10'b101110011;
	    10'b111001000: rot_addr = 10'b110010000;
	    10'b111001001: rot_addr = 10'b110010001;
	    10'b111001010: rot_addr = 10'b110101110;
	    10'b111001011: rot_addr = 10'b110101110;
	    10'b111001100: rot_addr = 10'b110101111;
	    10'b111001101: rot_addr = 10'b111001100;
	    10'b111001110: rot_addr = 10'b111001101;
	    10'b111001111: rot_addr = 10'b111001110;
	    10'b111010000: rot_addr = 10'b111101011;
	    10'b111010001: rot_addr = 10'b111101100;
	    10'b111010010: rot_addr = 10'b111101101;
	    10'b111010011: rot_addr = 10'b1000001010;
	    10'b111010100: rot_addr = 10'b1000001011;
	    10'b111010101: rot_addr = 10'b1000001100;
	    10'b111010110: rot_addr = 10'b1000101001;
	    10'b111010111: rot_addr = 10'b1000101010;
	    10'b111011000: rot_addr = 10'b1000101011;
	    10'b111011001: rot_addr = 10'b1001001000;
	    10'b111011010: rot_addr = 10'b1001001001;
	    10'b111011011: rot_addr = 10'b1001001010;
	    10'b111011100: rot_addr = 10'b0;
	    10'b111011101: rot_addr = 10'b101010001;
	    10'b111011110: rot_addr = 10'b101101110;
	    10'b111011111: rot_addr = 10'b101101111;
	    10'b111100000: rot_addr = 10'b101110000;
	    10'b111100001: rot_addr = 10'b110001101;
	    10'b111100010: rot_addr = 10'b110001101;
	    10'b111100011: rot_addr = 10'b110001110;
	    10'b111100100: rot_addr = 10'b110101011;
	    10'b111100101: rot_addr = 10'b110101100;
	    10'b111100110: rot_addr = 10'b110101101;
	    10'b111100111: rot_addr = 10'b111001010;
	    10'b111101000: rot_addr = 10'b111001011;
	    10'b111101001: rot_addr = 10'b111001100;
	    10'b111101010: rot_addr = 10'b111101001;
	    10'b111101011: rot_addr = 10'b111101010;
	    10'b111101100: rot_addr = 10'b1000000111;
	    10'b111101101: rot_addr = 10'b1000001000;
	    10'b111101110: rot_addr = 10'b1000001001;
	    10'b111101111: rot_addr = 10'b1000100110;
	    10'b111110000: rot_addr = 10'b1000100111;
	    10'b111110001: rot_addr = 10'b1000101000;
	    10'b111110010: rot_addr = 10'b1001000100;
	    10'b111110011: rot_addr = 10'b1001000101;
	    10'b111110100: rot_addr = 10'b1001000110;
	    10'b111110101: rot_addr = 10'b1001100011;
	    10'b111110110: rot_addr = 10'b1001100100;
	    10'b111110111: rot_addr = 10'b1001100101;
	    10'b111111000: rot_addr = 10'b0;
	    10'b111111001: rot_addr = 10'b0;
	    10'b111111010: rot_addr = 10'b110001001;
	    10'b111111011: rot_addr = 10'b110001010;
	    10'b111111100: rot_addr = 10'b110001011;
	    10'b111111101: rot_addr = 10'b110101000;
	    10'b111111110: rot_addr = 10'b110101001;
	    10'b111111111: rot_addr = 10'b110101010;
	    10'b1000000000: rot_addr = 10'b111000111;
	    10'b1000000001: rot_addr = 10'b111001000;
	    10'b1000000010: rot_addr = 10'b111001001;
	    10'b1000000011: rot_addr = 10'b111100110;
	    10'b1000000100: rot_addr = 10'b111100111;
	    10'b1000000101: rot_addr = 10'b111101000;
	    10'b1000000110: rot_addr = 10'b1000000101;
	    10'b1000000111: rot_addr = 10'b1000000110;
	    10'b1000001000: rot_addr = 10'b1000000111;
	    10'b1000001001: rot_addr = 10'b1000100011;
	    10'b1000001010: rot_addr = 10'b1000100100;
	    10'b1000001011: rot_addr = 10'b1000100101;
	    10'b1000001100: rot_addr = 10'b1001000010;
	    10'b1000001101: rot_addr = 10'b1001000011;
	    10'b1000001110: rot_addr = 10'b1001000100;
	    10'b1000001111: rot_addr = 10'b1001100001;
	    10'b1000010000: rot_addr = 10'b1001100010;
	    10'b1000010001: rot_addr = 10'b1001111111;
	    10'b1000010010: rot_addr = 10'b1010000000;
	    10'b1000010011: rot_addr = 10'b1010000001;
	    10'b1000010100: rot_addr = 10'b0;
	    10'b1000010101: rot_addr = 10'b0;
	    10'b1000010110: rot_addr = 10'b110100101;
	    10'b1000010111: rot_addr = 10'b110100110;
	    10'b1000011000: rot_addr = 10'b110100111;
	    10'b1000011001: rot_addr = 10'b111000100;
	    10'b1000011010: rot_addr = 10'b111000101;
	    10'b1000011011: rot_addr = 10'b111000110;
	    10'b1000011100: rot_addr = 10'b111100011;
	    10'b1000011101: rot_addr = 10'b111100100;
	    10'b1000011110: rot_addr = 10'b111100101;
	    10'b1000011111: rot_addr = 10'b1000000001;
	    10'b1000100000: rot_addr = 10'b1000000010;
	    10'b1000100001: rot_addr = 10'b1000000011;
	    10'b1000100010: rot_addr = 10'b1000100000;
	    10'b1000100011: rot_addr = 10'b1000100001;
	    10'b1000100100: rot_addr = 10'b1000100010;
	    10'b1000100101: rot_addr = 10'b1000111111;
	    10'b1000100110: rot_addr = 10'b1001000000;
	    10'b1000100111: rot_addr = 10'b1001000001;
	    10'b1000101000: rot_addr = 10'b1001011110;
	    10'b1000101001: rot_addr = 10'b1001011111;
	    10'b1000101010: rot_addr = 10'b1001100000;
	    10'b1000101011: rot_addr = 10'b1001111101;
	    10'b1000101100: rot_addr = 10'b1001111110;
	    10'b1000101101: rot_addr = 10'b1001111111;
	    10'b1000101110: rot_addr = 10'b1010011100;
	    10'b1000101111: rot_addr = 10'b1010011101;
	    10'b1000110000: rot_addr = 10'b0;
	    10'b1000110001: rot_addr = 10'b0;
	    10'b1000110010: rot_addr = 10'b111000001;
	    10'b1000110011: rot_addr = 10'b111000010;
	    10'b1000110100: rot_addr = 10'b111000011;
	    10'b1000110101: rot_addr = 10'b111011111;
	    10'b1000110110: rot_addr = 10'b111100000;
	    10'b1000110111: rot_addr = 10'b111100001;
	    10'b1000111000: rot_addr = 10'b111111110;
	    10'b1000111001: rot_addr = 10'b111111111;
	    10'b1000111010: rot_addr = 10'b1000000000;
	    10'b1000111011: rot_addr = 10'b1000011101;
	    10'b1000111100: rot_addr = 10'b1000011110;
	    10'b1000111101: rot_addr = 10'b1000011111;
	    10'b1000111110: rot_addr = 10'b1000111100;
	    10'b1000111111: rot_addr = 10'b1000111101;
	    10'b1001000000: rot_addr = 10'b1000111110;
	    10'b1001000001: rot_addr = 10'b1001011011;
	    10'b1001000010: rot_addr = 10'b1001011100;
	    10'b1001000011: rot_addr = 10'b1001011101;
	    10'b1001000100: rot_addr = 10'b1001111010;
	    10'b1001000101: rot_addr = 10'b1001111011;
	    10'b1001000110: rot_addr = 10'b1001111011;
	    10'b1001000111: rot_addr = 10'b1010011000;
	    10'b1001001000: rot_addr = 10'b1010011001;
	    10'b1001001001: rot_addr = 10'b1010011010;
	    10'b1001001010: rot_addr = 10'b1010110111;
	    10'b1001001011: rot_addr = 10'b1010111000;
	    10'b1001001100: rot_addr = 10'b0;
	    10'b1001001101: rot_addr = 10'b0;
	    10'b1001001110: rot_addr = 10'b0;
	    10'b1001001111: rot_addr = 10'b111011101;
	    10'b1001010000: rot_addr = 10'b111011110;
	    10'b1001010001: rot_addr = 10'b111011111;
	    10'b1001010010: rot_addr = 10'b111111100;
	    10'b1001010011: rot_addr = 10'b111111101;
	    10'b1001010100: rot_addr = 10'b1000011010;
	    10'b1001010101: rot_addr = 10'b1000011011;
	    10'b1001010110: rot_addr = 10'b1000011100;
	    10'b1001010111: rot_addr = 10'b1000111001;
	    10'b1001011000: rot_addr = 10'b1000111010;
	    10'b1001011001: rot_addr = 10'b1000111011;
	    10'b1001011010: rot_addr = 10'b1001011000;
	    10'b1001011011: rot_addr = 10'b1001011001;
	    10'b1001011100: rot_addr = 10'b1001011001;
	    10'b1001011101: rot_addr = 10'b1001110110;
	    10'b1001011110: rot_addr = 10'b1001110111;
	    10'b1001011111: rot_addr = 10'b1001111000;
	    10'b1001100000: rot_addr = 10'b1010010101;
	    10'b1001100001: rot_addr = 10'b1010010110;
	    10'b1001100010: rot_addr = 10'b1010010111;
	    10'b1001100011: rot_addr = 10'b1010110100;
	    10'b1001100100: rot_addr = 10'b1010110101;
	    10'b1001100101: rot_addr = 10'b1010110110;
	    10'b1001100110: rot_addr = 10'b1011010011;
	    10'b1001100111: rot_addr = 10'b1011010100;
	    10'b1001101000: rot_addr = 10'b0;
	    10'b1001101001: rot_addr = 10'b0;
	    10'b1001101010: rot_addr = 10'b0;
	    10'b1001101011: rot_addr = 10'b111111001;
	    10'b1001101100: rot_addr = 10'b111111010;
	    10'b1001101101: rot_addr = 10'b111111011;
	    10'b1001101110: rot_addr = 10'b1000011000;
	    10'b1001101111: rot_addr = 10'b1000011001;
	    10'b1001110000: rot_addr = 10'b1000011010;
	    10'b1001110001: rot_addr = 10'b1000110111;
	    10'b1001110010: rot_addr = 10'b1000111000;
	    10'b1001110011: rot_addr = 10'b1000111000;
	    10'b1001110100: rot_addr = 10'b1001010101;
	    10'b1001110101: rot_addr = 10'b1001010110;
	    10'b1001110110: rot_addr = 10'b1001110011;
	    10'b1001110111: rot_addr = 10'b1001110100;
	    10'b1001111000: rot_addr = 10'b1001110101;
	    10'b1001111001: rot_addr = 10'b1010010010;
	    10'b1001111010: rot_addr = 10'b1010010011;
	    10'b1001111011: rot_addr = 10'b1010010100;
	    10'b1001111100: rot_addr = 10'b1010110001;
	    10'b1001111101: rot_addr = 10'b1010110010;
	    10'b1001111110: rot_addr = 10'b1010110011;
	    10'b1001111111: rot_addr = 10'b1011010000;
	    10'b1010000000: rot_addr = 10'b1011010001;
	    10'b1010000001: rot_addr = 10'b1011010010;
	    10'b1010000010: rot_addr = 10'b1011101111;
	    10'b1010000011: rot_addr = 10'b1011101111;
	    10'b1010000100: rot_addr = 10'b0;
	    10'b1010000101: rot_addr = 10'b0;
	    10'b1010000110: rot_addr = 10'b0;
	    10'b1010000111: rot_addr = 10'b1000010101;
	    10'b1010001000: rot_addr = 10'b1000010110;
	    10'b1010001001: rot_addr = 10'b1000010110;
	    10'b1010001010: rot_addr = 10'b1000110011;
	    10'b1010001011: rot_addr = 10'b1000110100;
	    10'b1010001100: rot_addr = 10'b1000110101;
	    10'b1010001101: rot_addr = 10'b1001010010;
	    10'b1010001110: rot_addr = 10'b1001010011;
	    10'b1010001111: rot_addr = 10'b1001010100;
	    10'b1010010000: rot_addr = 10'b1001110001;
	    10'b1010010001: rot_addr = 10'b1001110010;
	    10'b1010010010: rot_addr = 10'b1001110011;
	    10'b1010010011: rot_addr = 10'b1010010000;
	    10'b1010010100: rot_addr = 10'b1010010001;
	    10'b1010010101: rot_addr = 10'b1010010010;
	    10'b1010010110: rot_addr = 10'b1010101111;
	    10'b1010010111: rot_addr = 10'b1010110000;
	    10'b1010011000: rot_addr = 10'b1011001101;
	    10'b1010011001: rot_addr = 10'b1011001101;
	    10'b1010011010: rot_addr = 10'b1011001110;
	    10'b1010011011: rot_addr = 10'b1011101011;
	    10'b1010011100: rot_addr = 10'b1011101100;
	    10'b1010011101: rot_addr = 10'b1011101101;
	    10'b1010011110: rot_addr = 10'b1100001010;
	    10'b1010011111: rot_addr = 10'b1100001011;
	    10'b1010100000: rot_addr = 10'b0;
	    10'b1010100001: rot_addr = 10'b0;
	    10'b1010100010: rot_addr = 10'b0;
	    10'b1010100011: rot_addr = 10'b0;
	    10'b1010100100: rot_addr = 10'b1000110001;
	    10'b1010100101: rot_addr = 10'b1000110010;
	    10'b1010100110: rot_addr = 10'b1001001111;
	    10'b1010100111: rot_addr = 10'b1001010000;
	    10'b1010101000: rot_addr = 10'b1001010001;
	    10'b1010101001: rot_addr = 10'b1001101110;
	    10'b1010101010: rot_addr = 10'b1001101111;
	    10'b1010101011: rot_addr = 10'b1001110000;
	    10'b1010101100: rot_addr = 10'b1010001101;
	    10'b1010101101: rot_addr = 10'b1010001110;
	    10'b1010101110: rot_addr = 10'b1010001111;
	    10'b1010101111: rot_addr = 10'b1010101100;
	    10'b1010110000: rot_addr = 10'b1010101100;
	    10'b1010110001: rot_addr = 10'b1010101101;
	    10'b1010110010: rot_addr = 10'b1011001010;
	    10'b1010110011: rot_addr = 10'b1011001011;
	    10'b1010110100: rot_addr = 10'b1011001100;
	    10'b1010110101: rot_addr = 10'b1011101001;
	    10'b1010110110: rot_addr = 10'b1011101010;
	    10'b1010110111: rot_addr = 10'b1011101011;
	    10'b1010111000: rot_addr = 10'b1100001000;
	    10'b1010111001: rot_addr = 10'b1100001001;
	    10'b1010111010: rot_addr = 10'b0;
	    10'b1010111011: rot_addr = 10'b0;
	    10'b1010111100: rot_addr = 10'b0;
	    10'b1010111101: rot_addr = 10'b0;
	    10'b1010111110: rot_addr = 10'b0;
	    10'b1010111111: rot_addr = 10'b0;
	    10'b1011000000: rot_addr = 10'b1001001101;
	    10'b1011000001: rot_addr = 10'b1001001110;
	    10'b1011000010: rot_addr = 10'b1001101011;
	    10'b1011000011: rot_addr = 10'b1001101100;
	    10'b1011000100: rot_addr = 10'b1001101101;
	    10'b1011000101: rot_addr = 10'b1010001010;
	    10'b1011000110: rot_addr = 10'b1010001010;
	    10'b1011000111: rot_addr = 10'b1010001011;
	    10'b1011001000: rot_addr = 10'b1010101000;
	    10'b1011001001: rot_addr = 10'b1010101001;
	    10'b1011001010: rot_addr = 10'b1010101010;
	    10'b1011001011: rot_addr = 10'b1011000111;
	    10'b1011001100: rot_addr = 10'b1011001000;
	    10'b1011001101: rot_addr = 10'b1011001001;
	    10'b1011001110: rot_addr = 10'b1011100110;
	    10'b1011001111: rot_addr = 10'b1011100111;
	    10'b1011010000: rot_addr = 10'b1011101000;
	    10'b1011010001: rot_addr = 10'b1100000101;
	    10'b1011010010: rot_addr = 10'b1100000110;
	    10'b1011010011: rot_addr = 10'b1100000111;
	    10'b1011010100: rot_addr = 10'b0;
	    10'b1011010101: rot_addr = 10'b0;
	    10'b1011010110: rot_addr = 10'b0;
	    10'b1011010111: rot_addr = 10'b0;
	    10'b1011011000: rot_addr = 10'b0;
	    10'b1011011001: rot_addr = 10'b0;
	    10'b1011011010: rot_addr = 10'b0;
	    10'b1011011011: rot_addr = 10'b0;
	    10'b1011011100: rot_addr = 10'b0;
	    10'b1011011101: rot_addr = 10'b1001101001;
	    10'b1011011110: rot_addr = 10'b1010000110;
	    10'b1011011111: rot_addr = 10'b1010000111;
	    10'b1011100000: rot_addr = 10'b1010001000;
	    10'b1011100001: rot_addr = 10'b1010100101;
	    10'b1011100010: rot_addr = 10'b1010100110;
	    10'b1011100011: rot_addr = 10'b1010100111;
	    10'b1011100100: rot_addr = 10'b1011000100;
	    10'b1011100101: rot_addr = 10'b1011000101;
	    10'b1011100110: rot_addr = 10'b1011000110;
	    10'b1011100111: rot_addr = 10'b1011100011;
	    10'b1011101000: rot_addr = 10'b1011100100;
	    10'b1011101001: rot_addr = 10'b1011100101;
	    10'b1011101010: rot_addr = 10'b1100000010;
	    10'b1011101011: rot_addr = 10'b1100000011;
	    10'b1011101100: rot_addr = 10'b1100000100;
	    10'b1011101101: rot_addr = 10'b0;
	    10'b1011101110: rot_addr = 10'b0;
	    10'b1011101111: rot_addr = 10'b0;
	    10'b1011110000: rot_addr = 10'b0;
	    10'b1011110001: rot_addr = 10'b0;
	    10'b1011110010: rot_addr = 10'b0;
	    10'b1011110011: rot_addr = 10'b0;
	    10'b1011110100: rot_addr = 10'b0;
	    10'b1011110101: rot_addr = 10'b0;
	    10'b1011110110: rot_addr = 10'b0;
	    10'b1011110111: rot_addr = 10'b0;
	    10'b1011111000: rot_addr = 10'b0;
	    10'b1011111001: rot_addr = 10'b1010000101;
	    10'b1011111010: rot_addr = 10'b1010000110;
	    10'b1011111011: rot_addr = 10'b1010100011;
	    10'b1011111100: rot_addr = 10'b1010100100;
	    10'b1011111101: rot_addr = 10'b1011000001;
	    10'b1011111110: rot_addr = 10'b1011000010;
	    10'b1011111111: rot_addr = 10'b1011000011;
	    10'b1100000000: rot_addr = 10'b1011100000;
	    10'b1100000001: rot_addr = 10'b1011100001;
	    10'b1100000010: rot_addr = 10'b1011100010;
	    10'b1100000011: rot_addr = 10'b1011111110;
	    10'b1100000100: rot_addr = 10'b1011111111;
	    10'b1100000101: rot_addr = 10'b1100000000;
	    10'b1100000110: rot_addr = 10'b0;
	    10'b1100000111: rot_addr = 10'b0;
	    10'b1100001000: rot_addr = 10'b0;
	    10'b1100001001: rot_addr = 10'b0;
	    10'b1100001010: rot_addr = 10'b0;
	    10'b1100001011: rot_addr = 10'b0;
	    10'b1100001100: rot_addr = 10'b0;
	    10'b1100001101: rot_addr = 10'b0;
	    10'b1100001110: rot_addr = 10'b0;
	    10'b1100001111: rot_addr = 10'b0;
	  endcase
	end 


endmodule
