

module BRAM_sim_biiiig (
    input  logic [31:0] address,
    output logic [31:0]  data_send,
    input logic clk,
    input logic reset
);
    logic [31:0] data;
    
    always_ff @(posedge clk)
    if (reset)
    data_send <= 32'd0;
    else
    data_send <= data;



    always_comb begin
        case (address)
            32'h00000000: data = 32'd0;
            32'h00000004: data = 32'd1;
            32'h00000008: data = 32'd2;
            32'h0000000C: data = 32'd3;
            32'h00000010: data = 32'd4;
            32'h00000014: data = 32'd5;
            32'h00000018: data = 32'd6;
            32'h0000001C: data = 32'd7;
            32'h00000020: data = 32'd8;
            32'h00000024: data = 32'd9;
            32'h00000028: data = 32'd10;
            32'h0000002C: data = 32'd11;
            32'h00000030: data = 32'd12;
            32'h00000034: data = 32'd13;
            32'h00000038: data = 32'd14;
            32'h0000003C: data = 32'd15;
            32'h00000040: data = 32'd16;
            32'h00000044: data = 32'd17;
            32'h00000048: data = 32'd18;
            32'h0000004C: data = 32'd19;
            32'h00000050: data = 32'd20;
            32'h00000054: data = 32'd21;
            32'h00000058: data = 32'd22;
            32'h0000005C: data = 32'd23;
            32'h00000060: data = 32'd24;
            32'h00000064: data = 32'd25;
            32'h00000068: data = 32'd26;
            32'h0000006C: data = 32'd27;
            32'h00000070: data = 32'd28;
            32'h00000074: data = 32'd29;
            32'h00000078: data = 32'd30;
            32'h0000007C: data = 32'd31;
            32'h00000080: data = 32'd32;
            32'h00000084: data = 32'd33;
            32'h00000088: data = 32'd34;
            32'h0000008C: data = 32'd35;
            32'h00000090: data = 32'd36;
            32'h00000094: data = 32'd37;
            32'h00000098: data = 32'd38;
            32'h0000009C: data = 32'd39;
            32'h000000A0: data = 32'd40;
            32'h000000A4: data = 32'd41;
            32'h000000A8: data = 32'd42;
            32'h000000AC: data = 32'd43;
            32'h000000B0: data = 32'd44;
            32'h000000B4: data = 32'd45;
            32'h000000B8: data = 32'd46;
            32'h000000BC: data = 32'd47;
            32'h000000C0: data = 32'd48;
            32'h000000C4: data = 32'd49;
            32'h000000C8: data = 32'd50;
            32'h000000CC: data = 32'd51;
            32'h000000D0: data = 32'd52;
            32'h000000D4: data = 32'd53;
            32'h000000D8: data = 32'd54;
            32'h000000DC: data = 32'd55;
            32'h000000E0: data = 32'd56;
            32'h000000E4: data = 32'd57;
            32'h000000E8: data = 32'd58;
            32'h000000EC: data = 32'd59;
            32'h000000F0: data = 32'd60;
            32'h000000F4: data = 32'd61;
            32'h000000F8: data = 32'd62;
            32'h000000FC: data = 32'd63;
            32'h00000100: data = 32'd64;
            32'h00000104: data = 32'd65;
            32'h00000108: data = 32'd66;
            32'h0000010C: data = 32'd67;
            32'h00000110: data = 32'd68;
            32'h00000114: data = 32'd69;
            32'h00000118: data = 32'd70;
            32'h0000011C: data = 32'd71;
            32'h00000120: data = 32'd72;
            32'h00000124: data = 32'd73;
            32'h00000128: data = 32'd74;
            32'h0000012C: data = 32'd75;
            32'h00000130: data = 32'd76;
            32'h00000134: data = 32'd77;
            32'h00000138: data = 32'd78;
            32'h0000013C: data = 32'd79;
            32'h00000140: data = 32'd80;
            32'h00000144: data = 32'd81;
            32'h00000148: data = 32'd82;
            32'h0000014C: data = 32'd83;
            32'h00000150: data = 32'd84;
            32'h00000154: data = 32'd85;
            32'h00000158: data = 32'd86;
            32'h0000015C: data = 32'd87;
            32'h00000160: data = 32'd88;
            32'h00000164: data = 32'd89;
            32'h00000168: data = 32'd90;
            32'h0000016C: data = 32'd91;
            32'h00000170: data = 32'd92;
            32'h00000174: data = 32'd93;
            32'h00000178: data = 32'd94;
            32'h0000017C: data = 32'd95;
            32'h00000180: data = 32'd96;
            32'h00000184: data = 32'd97;
            32'h00000188: data = 32'd98;
            32'h0000018C: data = 32'd99;
            32'h00000190: data = 32'd100;
            32'h00000194: data = 32'd101;
            32'h00000198: data = 32'd102;
            32'h0000019C: data = 32'd103;
            32'h000001A0: data = 32'd104;
            32'h000001A4: data = 32'd105;
            32'h000001A8: data = 32'd106;
            32'h000001AC: data = 32'd107;
            32'h000001B0: data = 32'd108;
            32'h000001B4: data = 32'd109;
            32'h000001B8: data = 32'd110;
            32'h000001BC: data = 32'd111;
            32'h000001C0: data = 32'd112;
            32'h000001C4: data = 32'd113;
            32'h000001C8: data = 32'd114;
            32'h000001CC: data = 32'd115;
            32'h000001D0: data = 32'd116;
            32'h000001D4: data = 32'd117;
            32'h000001D8: data = 32'd118;
            32'h000001DC: data = 32'd119;
            32'h000001E0: data = 32'd120;
            32'h000001E4: data = 32'd121;
            32'h000001E8: data = 32'd122;
            32'h000001EC: data = 32'd123;
            32'h000001F0: data = 32'd124;
            32'h000001F4: data = 32'd125;
            32'h000001F8: data = 32'd126;
            32'h000001FC: data = 32'd127;
            32'h00000200: data = 32'd128;
            32'h00000204: data = 32'd129;
            32'h00000208: data = 32'd130;
            32'h0000020C: data = 32'd131;
            32'h00000210: data = 32'd132;
            32'h00000214: data = 32'd133;
            32'h00000218: data = 32'd134;
            32'h0000021C: data = 32'd135;
            32'h00000220: data = 32'd136;
            32'h00000224: data = 32'd137;
            32'h00000228: data = 32'd138;
            32'h0000022C: data = 32'd139;
            32'h00000230: data = 32'd140;
            32'h00000234: data = 32'd141;
            32'h00000238: data = 32'd142;
            32'h0000023C: data = 32'd143;
            32'h00000240: data = 32'd144;
            32'h00000244: data = 32'd145;
            32'h00000248: data = 32'd146;
            32'h0000024C: data = 32'd147;
            32'h00000250: data = 32'd148;
            32'h00000254: data = 32'd149;
            32'h00000258: data = 32'd150;
            32'h0000025C: data = 32'd151;
            32'h00000260: data = 32'd152;
            32'h00000264: data = 32'd153;
            32'h00000268: data = 32'd154;
            32'h0000026C: data = 32'd155;
            32'h00000270: data = 32'd156;
            32'h00000274: data = 32'd157;
            32'h00000278: data = 32'd158;
            32'h0000027C: data = 32'd159;
            32'h00000280: data = 32'd160;
            32'h00000284: data = 32'd161;
            32'h00000288: data = 32'd162;
            32'h0000028C: data = 32'd163;
            32'h00000290: data = 32'd164;
            32'h00000294: data = 32'd165;
            32'h00000298: data = 32'd166;
            32'h0000029C: data = 32'd167;
            32'h000002A0: data = 32'd168;
            32'h000002A4: data = 32'd169;
            32'h000002A8: data = 32'd170;
            32'h000002AC: data = 32'd171;
            32'h000002B0: data = 32'd172;
            32'h000002B4: data = 32'd173;
            32'h000002B8: data = 32'd174;
            32'h000002BC: data = 32'd175;
            32'h000002C0: data = 32'd176;
            32'h000002C4: data = 32'd177;
            32'h000002C8: data = 32'd178;
            32'h000002CC: data = 32'd179;
            32'h000002D0: data = 32'd180;
            32'h000002D4: data = 32'd181;
            32'h000002D8: data = 32'd182;
            32'h000002DC: data = 32'd183;
            32'h000002E0: data = 32'd184;
            32'h000002E4: data = 32'd185;
            32'h000002E8: data = 32'd186;
            32'h000002EC: data = 32'd187;
            32'h000002F0: data = 32'd188;
            32'h000002F4: data = 32'd189;
            32'h000002F8: data = 32'd190;
            32'h000002FC: data = 32'd191;
            32'h00000300: data = 32'd192;
            32'h00000304: data = 32'd193;
            32'h00000308: data = 32'd194;
            32'h0000030C: data = 32'd195;
            32'h00000310: data = 32'd196;
            32'h00000314: data = 32'd197;
            32'h00000318: data = 32'd198;
            32'h0000031C: data = 32'd199;
            32'h00000320: data = 32'd200;
            32'h00000324: data = 32'd201;
            32'h00000328: data = 32'd202;
            32'h0000032C: data = 32'd203;
            32'h00000330: data = 32'd204;
            32'h00000334: data = 32'd205;
            32'h00000338: data = 32'd206;
            32'h0000033C: data = 32'd207;
            32'h00000340: data = 32'd208;
            32'h00000344: data = 32'd209;
            32'h00000348: data = 32'd210;
            32'h0000034C: data = 32'd211;
            32'h00000350: data = 32'd212;
            32'h00000354: data = 32'd213;
            32'h00000358: data = 32'd214;
            32'h0000035C: data = 32'd215;
            32'h00000360: data = 32'd216;
            32'h00000364: data = 32'd217;
            32'h00000368: data = 32'd218;
            32'h0000036C: data = 32'd219;
            32'h00000370: data = 32'd220;
            32'h00000374: data = 32'd221;
            32'h00000378: data = 32'd222;
            32'h0000037C: data = 32'd223;
            32'h00000380: data = 32'd224;
            32'h00000384: data = 32'd225;
            32'h00000388: data = 32'd226;
            32'h0000038C: data = 32'd227;
            32'h00000390: data = 32'd228;
            32'h00000394: data = 32'd229;
            32'h00000398: data = 32'd230;
            32'h0000039C: data = 32'd231;
            32'h000003A0: data = 32'd232;
            32'h000003A4: data = 32'd233;
            32'h000003A8: data = 32'd234;
            32'h000003AC: data = 32'd235;
            32'h000003B0: data = 32'd236;
            32'h000003B4: data = 32'd237;
            32'h000003B8: data = 32'd238;
            32'h000003BC: data = 32'd239;
            32'h000003C0: data = 32'd240;
            32'h000003C4: data = 32'd241;
            32'h000003C8: data = 32'd242;
            32'h000003CC: data = 32'd243;
            32'h000003D0: data = 32'd244;
            32'h000003D4: data = 32'd245;
            32'h000003D8: data = 32'd246;
            32'h000003DC: data = 32'd247;
            32'h000003E0: data = 32'd248;
            32'h000003E4: data = 32'd249;
            32'h000003E8: data = 32'd250;
            32'h000003EC: data = 32'd251;
            32'h000003F0: data = 32'd252;
            32'h000003F4: data = 32'd253;
            32'h000003F8: data = 32'd254;
            32'h000003FC: data = 32'd255;
            32'h00000400: data = 32'd0;
            32'h00000404: data = 32'd1;
            32'h00000408: data = 32'd2;
            32'h0000040C: data = 32'd3;
            32'h00000410: data = 32'd4;
            32'h00000414: data = 32'd5;
            32'h00000418: data = 32'd6;
            32'h0000041C: data = 32'd7;
            32'h00000420: data = 32'd8;
            32'h00000424: data = 32'd9;
            32'h00000428: data = 32'd10;
            32'h0000042C: data = 32'd11;
            32'h00000430: data = 32'd12;
            32'h00000434: data = 32'd13;
            32'h00000438: data = 32'd14;
            32'h0000043C: data = 32'd15;
            32'h00000440: data = 32'd16;
            32'h00000444: data = 32'd17;
            32'h00000448: data = 32'd18;
            32'h0000044C: data = 32'd19;
            32'h00000450: data = 32'd20;
            32'h00000454: data = 32'd21;
            32'h00000458: data = 32'd22;
            32'h0000045C: data = 32'd23;
            32'h00000460: data = 32'd24;
            32'h00000464: data = 32'd25;
            32'h00000468: data = 32'd26;
            32'h0000046C: data = 32'd27;
            32'h00000470: data = 32'd28;
            32'h00000474: data = 32'd29;
            32'h00000478: data = 32'd30;
            32'h0000047C: data = 32'd31;
            32'h00000480: data = 32'd32;
            32'h00000484: data = 32'd33;
            32'h00000488: data = 32'd34;
            32'h0000048C: data = 32'd35;
            32'h00000490: data = 32'd36;
            32'h00000494: data = 32'd37;
            32'h00000498: data = 32'd38;
            32'h0000049C: data = 32'd39;
            32'h000004A0: data = 32'd40;
            32'h000004A4: data = 32'd41;
            32'h000004A8: data = 32'd42;
            32'h000004AC: data = 32'd43;
            32'h000004B0: data = 32'd44;
            32'h000004B4: data = 32'd45;
            32'h000004B8: data = 32'd46;
            32'h000004BC: data = 32'd47;
            32'h000004C0: data = 32'd48;
            32'h000004C4: data = 32'd49;
            32'h000004C8: data = 32'd50;
            32'h000004CC: data = 32'd51;
            32'h000004D0: data = 32'd52;
            32'h000004D4: data = 32'd53;
            32'h000004D8: data = 32'd54;
            32'h000004DC: data = 32'd55;
            32'h000004E0: data = 32'd56;
            32'h000004E4: data = 32'd57;
            32'h000004E8: data = 32'd58;
            32'h000004EC: data = 32'd59;
            32'h000004F0: data = 32'd60;
            32'h000004F4: data = 32'd61;
            32'h000004F8: data = 32'd62;
            32'h000004FC: data = 32'd63;
            32'h00000500: data = 32'd64;
            32'h00000504: data = 32'd65;
            32'h00000508: data = 32'd66;
            32'h0000050C: data = 32'd67;
            32'h00000510: data = 32'd68;
            32'h00000514: data = 32'd69;
            32'h00000518: data = 32'd70;
            32'h0000051C: data = 32'd71;
            32'h00000520: data = 32'd72;
            32'h00000524: data = 32'd73;
            32'h00000528: data = 32'd74;
            32'h0000052C: data = 32'd75;
            32'h00000530: data = 32'd76;
            32'h00000534: data = 32'd77;
            32'h00000538: data = 32'd78;
            32'h0000053C: data = 32'd79;
            32'h00000540: data = 32'd80;
            32'h00000544: data = 32'd81;
            32'h00000548: data = 32'd82;
            32'h0000054C: data = 32'd83;
            32'h00000550: data = 32'd84;
            32'h00000554: data = 32'd85;
            32'h00000558: data = 32'd86;
            32'h0000055C: data = 32'd87;
            32'h00000560: data = 32'd88;
            32'h00000564: data = 32'd89;
            32'h00000568: data = 32'd90;
            32'h0000056C: data = 32'd91;
            32'h00000570: data = 32'd92;
            32'h00000574: data = 32'd93;
            32'h00000578: data = 32'd94;
            32'h0000057C: data = 32'd95;
            32'h00000580: data = 32'd96;
            32'h00000584: data = 32'd97;
            32'h00000588: data = 32'd98;
            32'h0000058C: data = 32'd99;
            32'h00000590: data = 32'd100;
            32'h00000594: data = 32'd101;
            32'h00000598: data = 32'd102;
            32'h0000059C: data = 32'd103;
            32'h000005A0: data = 32'd104;
            32'h000005A4: data = 32'd105;
            32'h000005A8: data = 32'd106;
            32'h000005AC: data = 32'd107;
            32'h000005B0: data = 32'd108;
            32'h000005B4: data = 32'd109;
            32'h000005B8: data = 32'd110;
            32'h000005BC: data = 32'd111;
            32'h000005C0: data = 32'd112;
            32'h000005C4: data = 32'd113;
            32'h000005C8: data = 32'd114;
            32'h000005CC: data = 32'd115;
            32'h000005D0: data = 32'd116;
            32'h000005D4: data = 32'd117;
            32'h000005D8: data = 32'd118;
            32'h000005DC: data = 32'd119;
            32'h000005E0: data = 32'd120;
            32'h000005E4: data = 32'd121;
            32'h000005E8: data = 32'd122;
            32'h000005EC: data = 32'd123;
            32'h000005F0: data = 32'd124;
            32'h000005F4: data = 32'd125;
            32'h000005F8: data = 32'd126;
            32'h000005FC: data = 32'd127;
            32'h00000600: data = 32'd128;
            32'h00000604: data = 32'd129;
            32'h00000608: data = 32'd130;
            32'h0000060C: data = 32'd131;
            32'h00000610: data = 32'd132;
            32'h00000614: data = 32'd133;
            32'h00000618: data = 32'd134;
            32'h0000061C: data = 32'd135;
            32'h00000620: data = 32'd136;
            32'h00000624: data = 32'd137;
            32'h00000628: data = 32'd138;
            32'h0000062C: data = 32'd139;
            32'h00000630: data = 32'd140;
            32'h00000634: data = 32'd141;
            32'h00000638: data = 32'd142;
            32'h0000063C: data = 32'd143;
            32'h00000640: data = 32'd144;
            32'h00000644: data = 32'd145;
            32'h00000648: data = 32'd146;
            32'h0000064C: data = 32'd147;
            32'h00000650: data = 32'd148;
            32'h00000654: data = 32'd149;
            32'h00000658: data = 32'd150;
            32'h0000065C: data = 32'd151;
            32'h00000660: data = 32'd152;
            32'h00000664: data = 32'd153;
            32'h00000668: data = 32'd154;
            32'h0000066C: data = 32'd155;
            32'h00000670: data = 32'd156;
            32'h00000674: data = 32'd157;
            32'h00000678: data = 32'd158;
            32'h0000067C: data = 32'd159;
            32'h00000680: data = 32'd160;
            32'h00000684: data = 32'd161;
            32'h00000688: data = 32'd162;
            32'h0000068C: data = 32'd163;
            32'h00000690: data = 32'd164;
            32'h00000694: data = 32'd165;
            32'h00000698: data = 32'd166;
            32'h0000069C: data = 32'd167;
            32'h000006A0: data = 32'd168;
            32'h000006A4: data = 32'd169;
            32'h000006A8: data = 32'd170;
            32'h000006AC: data = 32'd171;
            32'h000006B0: data = 32'd172;
            32'h000006B4: data = 32'd173;
            32'h000006B8: data = 32'd174;
            32'h000006BC: data = 32'd175;
            32'h000006C0: data = 32'd176;
            32'h000006C4: data = 32'd177;
            32'h000006C8: data = 32'd178;
            32'h000006CC: data = 32'd179;
            32'h000006D0: data = 32'd180;
            32'h000006D4: data = 32'd181;
            32'h000006D8: data = 32'd182;
            32'h000006DC: data = 32'd183;
            32'h000006E0: data = 32'd184;
            32'h000006E4: data = 32'd185;
            32'h000006E8: data = 32'd186;
            32'h000006EC: data = 32'd187;
            32'h000006F0: data = 32'd188;
            32'h000006F4: data = 32'd189;
            32'h000006F8: data = 32'd190;
            32'h000006FC: data = 32'd191;
            32'h00000700: data = 32'd192;
            32'h00000704: data = 32'd193;
            32'h00000708: data = 32'd194;
            32'h0000070C: data = 32'd195;
            32'h00000710: data = 32'd196;
            32'h00000714: data = 32'd197;
            32'h00000718: data = 32'd198;
            32'h0000071C: data = 32'd199;
            32'h00000720: data = 32'd200;
            32'h00000724: data = 32'd201;
            32'h00000728: data = 32'd202;
            32'h0000072C: data = 32'd203;
            32'h00000730: data = 32'd204;
            32'h00000734: data = 32'd205;
            32'h00000738: data = 32'd206;
            32'h0000073C: data = 32'd207;
            32'h00000740: data = 32'd208;
            32'h00000744: data = 32'd209;
            32'h00000748: data = 32'd210;
            32'h0000074C: data = 32'd211;
            32'h00000750: data = 32'd212;
            32'h00000754: data = 32'd213;
            32'h00000758: data = 32'd214;
            32'h0000075C: data = 32'd215;
            32'h00000760: data = 32'd216;
            32'h00000764: data = 32'd217;
            32'h00000768: data = 32'd218;
            32'h0000076C: data = 32'd219;
            32'h00000770: data = 32'd220;
            32'h00000774: data = 32'd221;
            32'h00000778: data = 32'd222;
            32'h0000077C: data = 32'd223;
            32'h00000780: data = 32'd224;
            32'h00000784: data = 32'd225;
            32'h00000788: data = 32'd226;
            32'h0000078C: data = 32'd227;
            32'h00000790: data = 32'd228;
            32'h00000794: data = 32'd229;
            32'h00000798: data = 32'd230;
            32'h0000079C: data = 32'd231;
            32'h000007A0: data = 32'd232;
            32'h000007A4: data = 32'd233;
            32'h000007A8: data = 32'd234;
            32'h000007AC: data = 32'd235;
            32'h000007B0: data = 32'd236;
            32'h000007B4: data = 32'd237;
            32'h000007B8: data = 32'd238;
            32'h000007BC: data = 32'd239;
            32'h000007C0: data = 32'd240;
            32'h000007C4: data = 32'd241;
            32'h000007C8: data = 32'd242;
            32'h000007CC: data = 32'd243;
            32'h000007D0: data = 32'd244;
            32'h000007D4: data = 32'd245;
            32'h000007D8: data = 32'd246;
            32'h000007DC: data = 32'd247;
            32'h000007E0: data = 32'd248;
            32'h000007E4: data = 32'd249;
            32'h000007E8: data = 32'd250;
            32'h000007EC: data = 32'd251;
            32'h000007F0: data = 32'd252;
            32'h000007F4: data = 32'd253;
            32'h000007F8: data = 32'd254;
            32'h000007FC: data = 32'd255;
            32'h00000800: data = 32'd0;
            32'h00000804: data = 32'd1;
            32'h00000808: data = 32'd2;
            32'h0000080C: data = 32'd3;
            32'h00000810: data = 32'd4;
            32'h00000814: data = 32'd5;
            32'h00000818: data = 32'd6;
            32'h0000081C: data = 32'd7;
            32'h00000820: data = 32'd8;
            32'h00000824: data = 32'd9;
            32'h00000828: data = 32'd10;
            32'h0000082C: data = 32'd11;
            32'h00000830: data = 32'd12;
            32'h00000834: data = 32'd13;
            32'h00000838: data = 32'd14;
            32'h0000083C: data = 32'd15;
            32'h00000840: data = 32'd16;
            32'h00000844: data = 32'd17;
            32'h00000848: data = 32'd18;
            32'h0000084C: data = 32'd19;
            32'h00000850: data = 32'd20;
            32'h00000854: data = 32'd21;
            32'h00000858: data = 32'd22;
            32'h0000085C: data = 32'd23;
            32'h00000860: data = 32'd24;
            32'h00000864: data = 32'd25;
            32'h00000868: data = 32'd26;
            32'h0000086C: data = 32'd27;
            32'h00000870: data = 32'd28;
            32'h00000874: data = 32'd29;
            32'h00000878: data = 32'd30;
            32'h0000087C: data = 32'd31;
            32'h00000880: data = 32'd32;
            32'h00000884: data = 32'd33;
            32'h00000888: data = 32'd34;
            32'h0000088C: data = 32'd35;
            32'h00000890: data = 32'd36;
            32'h00000894: data = 32'd37;
            32'h00000898: data = 32'd38;
            32'h0000089C: data = 32'd39;
            32'h000008A0: data = 32'd40;
            32'h000008A4: data = 32'd41;
            32'h000008A8: data = 32'd42;
            32'h000008AC: data = 32'd43;
            32'h000008B0: data = 32'd44;
            32'h000008B4: data = 32'd45;
            32'h000008B8: data = 32'd46;
            32'h000008BC: data = 32'd47;
            32'h000008C0: data = 32'd48;
            32'h000008C4: data = 32'd49;
            32'h000008C8: data = 32'd50;
            32'h000008CC: data = 32'd51;
            32'h000008D0: data = 32'd52;
            32'h000008D4: data = 32'd53;
            32'h000008D8: data = 32'd54;
            32'h000008DC: data = 32'd55;
            32'h000008E0: data = 32'd56;
            32'h000008E4: data = 32'd57;
            32'h000008E8: data = 32'd58;
            32'h000008EC: data = 32'd59;
            32'h000008F0: data = 32'd60;
            32'h000008F4: data = 32'd61;
            32'h000008F8: data = 32'd62;
            32'h000008FC: data = 32'd63;
            32'h00000900: data = 32'd64;
            32'h00000904: data = 32'd65;
            32'h00000908: data = 32'd66;
            32'h0000090C: data = 32'd67;
            32'h00000910: data = 32'd68;
            32'h00000914: data = 32'd69;
            32'h00000918: data = 32'd70;
            32'h0000091C: data = 32'd71;
            32'h00000920: data = 32'd72;
            32'h00000924: data = 32'd73;
            32'h00000928: data = 32'd74;
            32'h0000092C: data = 32'd75;
            32'h00000930: data = 32'd76;
            32'h00000934: data = 32'd77;
            32'h00000938: data = 32'd78;
            32'h0000093C: data = 32'd79;
            32'h00000940: data = 32'd80;
            32'h00000944: data = 32'd81;
            32'h00000948: data = 32'd82;
            32'h0000094C: data = 32'd83;
            32'h00000950: data = 32'd84;
            32'h00000954: data = 32'd85;
            32'h00000958: data = 32'd86;
            32'h0000095C: data = 32'd87;
            32'h00000960: data = 32'd88;
            32'h00000964: data = 32'd89;
            32'h00000968: data = 32'd90;
            32'h0000096C: data = 32'd91;
            32'h00000970: data = 32'd92;
            32'h00000974: data = 32'd93;
            32'h00000978: data = 32'd94;
            32'h0000097C: data = 32'd95;
            32'h00000980: data = 32'd96;
            32'h00000984: data = 32'd97;
            32'h00000988: data = 32'd98;
            32'h0000098C: data = 32'd99;
            32'h00000990: data = 32'd100;
            32'h00000994: data = 32'd101;
            32'h00000998: data = 32'd102;
            32'h0000099C: data = 32'd103;
            32'h000009A0: data = 32'd104;
            32'h000009A4: data = 32'd105;
            32'h000009A8: data = 32'd106;
            32'h000009AC: data = 32'd107;
            32'h000009B0: data = 32'd108;
            32'h000009B4: data = 32'd109;
            32'h000009B8: data = 32'd110;
            32'h000009BC: data = 32'd111;
            32'h000009C0: data = 32'd112;
            32'h000009C4: data = 32'd113;
            32'h000009C8: data = 32'd114;
            32'h000009CC: data = 32'd115;
            32'h000009D0: data = 32'd116;
            32'h000009D4: data = 32'd117;
            32'h000009D8: data = 32'd118;
            32'h000009DC: data = 32'd119;
            32'h000009E0: data = 32'd120;
            32'h000009E4: data = 32'd121;
            32'h000009E8: data = 32'd122;
            32'h000009EC: data = 32'd123;
            32'h000009F0: data = 32'd124;
            32'h000009F4: data = 32'd125;
            32'h000009F8: data = 32'd126;
            32'h000009FC: data = 32'd127;
            32'h00000A00: data = 32'd128;
            32'h00000A04: data = 32'd129;
            32'h00000A08: data = 32'd130;
            32'h00000A0C: data = 32'd131;
            32'h00000A10: data = 32'd132;
            32'h00000A14: data = 32'd133;
            32'h00000A18: data = 32'd134;
            32'h00000A1C: data = 32'd135;
            32'h00000A20: data = 32'd136;
            32'h00000A24: data = 32'd137;
            32'h00000A28: data = 32'd138;
            32'h00000A2C: data = 32'd139;
            32'h00000A30: data = 32'd140;
            32'h00000A34: data = 32'd141;
            32'h00000A38: data = 32'd142;
            32'h00000A3C: data = 32'd143;
            32'h00000A40: data = 32'd144;
            32'h00000A44: data = 32'd145;
            32'h00000A48: data = 32'd146;
            32'h00000A4C: data = 32'd147;
            32'h00000A50: data = 32'd148;
            32'h00000A54: data = 32'd149;
            32'h00000A58: data = 32'd150;
            32'h00000A5C: data = 32'd151;
            32'h00000A60: data = 32'd152;
            32'h00000A64: data = 32'd153;
            32'h00000A68: data = 32'd154;
            32'h00000A6C: data = 32'd155;
            32'h00000A70: data = 32'd156;
            32'h00000A74: data = 32'd157;
            32'h00000A78: data = 32'd158;
            32'h00000A7C: data = 32'd159;
            32'h00000A80: data = 32'd160;
            32'h00000A84: data = 32'd161;
            32'h00000A88: data = 32'd162;
            32'h00000A8C: data = 32'd163;
            32'h00000A90: data = 32'd164;
            32'h00000A94: data = 32'd165;
            32'h00000A98: data = 32'd166;
            32'h00000A9C: data = 32'd167;
            32'h00000AA0: data = 32'd168;
            32'h00000AA4: data = 32'd169;
            32'h00000AA8: data = 32'd170;
            32'h00000AAC: data = 32'd171;
            32'h00000AB0: data = 32'd172;
            32'h00000AB4: data = 32'd173;
            32'h00000AB8: data = 32'd174;
            32'h00000ABC: data = 32'd175;
            32'h00000AC0: data = 32'd176;
            32'h00000AC4: data = 32'd177;
            32'h00000AC8: data = 32'd178;
            32'h00000ACC: data = 32'd179;
            32'h00000AD0: data = 32'd180;
            32'h00000AD4: data = 32'd181;
            32'h00000AD8: data = 32'd182;
            32'h00000ADC: data = 32'd183;
            32'h00000AE0: data = 32'd184;
            32'h00000AE4: data = 32'd185;
            32'h00000AE8: data = 32'd186;
            32'h00000AEC: data = 32'd187;
            32'h00000AF0: data = 32'd188;
            32'h00000AF4: data = 32'd189;
            32'h00000AF8: data = 32'd190;
            32'h00000AFC: data = 32'd191;
            32'h0000B000: data = 32'd192;
            32'h0000B004: data = 32'd193;
            32'h0000B008: data = 32'd194;
            32'h0000B00C: data = 32'd195;
            32'h00000B10: data = 32'd196;
            32'h00000B14: data = 32'd197;
            32'h00000B18: data = 32'd198;
            32'h00000B1C: data = 32'd199;
            32'h00000B20: data = 32'd200;
            32'h00000B24: data = 32'd201;
            32'h00000B28: data = 32'd202;
            32'h00000B2C: data = 32'd203;
            32'h00000B30: data = 32'd204;
            32'h00000B34: data = 32'd205;
            32'h00000B38: data = 32'd206;
            32'h00000B3C: data = 32'd207;
            32'h00000B40: data = 32'd208;
            32'h00000B44: data = 32'd209;
            32'h00000B48: data = 32'd210;
            32'h00000B4C: data = 32'd211;
            32'h00000B50: data = 32'd212;
            32'h00000B54: data = 32'd213;
            32'h00000B58: data = 32'd214;
            32'h00000B5C: data = 32'd215;
            32'h00000B60: data = 32'd216;
            32'h00000B64: data = 32'd217;
            32'h00000B68: data = 32'd218;
            32'h00000B6C: data = 32'd219;
            32'h00000B70: data = 32'd220;
            32'h00000B74: data = 32'd221;
            32'h00000B78: data = 32'd222;
            32'h00000B7C: data = 32'd223;
            32'h00000B80: data = 32'd224;
            32'h00000B84: data = 32'd225;
            32'h00000B88: data = 32'd226;
            32'h00000B8C: data = 32'd227;
            32'h00000B90: data = 32'd228;
            32'h00000B94: data = 32'd229;
            32'h00000B98: data = 32'd230;
            32'h00000B9C: data = 32'd231;
            32'h00000BA0: data = 32'd232;
            32'h00000BA4: data = 32'd233;
            32'h00000BA8: data = 32'd234;
            32'h00000BAC: data = 32'd235;
            32'h00000B00: data = 32'd236;
            32'h00000BB4: data = 32'd237;
            32'h00000BB8: data = 32'd238;
            32'h00000BBC: data = 32'd239;
            32'h00000BC0: data = 32'd240;
            32'h00000BC4: data = 32'd241;
            32'h00000BC8: data = 32'd242;
            32'h00000BCC: data = 32'd243;
            32'h00000BD0: data = 32'd244;
            32'h00000BD4: data = 32'd245;
            32'h00000BD8: data = 32'd246;
            32'h00000BDC: data = 32'd247;
            32'h00000BE0: data = 32'd248;
            32'h00000BE4: data = 32'd249;
            32'h00000BE8: data = 32'd250;
            32'h00000BEC: data = 32'd251;
            32'h00000BF0: data = 32'd252;
            32'h00000BF4: data = 32'd253;
            32'h00000BF8: data = 32'd254;
            32'h00000BFC: data = 32'd255;
            32'h00000C00: data = 32'd0;
            32'h00000C04: data = 32'd1;
            32'h00000C08: data = 32'd2;
            32'h00000C0C: data = 32'd3;
            32'h00000C10: data = 32'd4;
            32'h00000C14: data = 32'd5;
            32'h00000C18: data = 32'd6;
            32'h00000C1C: data = 32'd7;
            32'h00000C20: data = 32'd8;
            32'h00000C24: data = 32'd9;
            32'h00000C28: data = 32'd10;
            32'h00000C2C: data = 32'd11;
            32'h00000C30: data = 32'd12;
            32'h00000C34: data = 32'd13;
            32'h00000C38: data = 32'd14;
            32'h00000C3C: data = 32'd15;
            32'h00000C40: data = 32'd16;
            32'h00000C44: data = 32'd17;
            32'h00000C48: data = 32'd18;
            32'h00000C4C: data = 32'd19;
            32'h00000C50: data = 32'd20;
            32'h00000C54: data = 32'd21;
            32'h00000C58: data = 32'd22;
            32'h00000C5C: data = 32'd23;
            32'h00000C60: data = 32'd24;
            32'h00000C64: data = 32'd25;
            32'h00000C68: data = 32'd26;
            32'h00000C6C: data = 32'd27;
            32'h00000C70: data = 32'd28;
            32'h00000C74: data = 32'd29;
            32'h00000C78: data = 32'd30;
            32'h00000C7C: data = 32'd31;
            32'h00000C80: data = 32'd32;
            32'h00000C84: data = 32'd33;
            32'h00000C88: data = 32'd34;
            32'h00000C8C: data = 32'd35;
            32'h00000C90: data = 32'd36;
            32'h00000C94: data = 32'd37;
            32'h00000C98: data = 32'd38;
            32'h00000C9C: data = 32'd39;
            32'h00000CA0: data = 32'd40;
            32'h00000CA4: data = 32'd41;
            32'h00000CA8: data = 32'd42;
            32'h00000CAC: data = 32'd43;
            32'h00000CB0: data = 32'd44;
            32'h00000CB4: data = 32'd45;
            32'h00000CB8: data = 32'd46;
            32'h00000CBC: data = 32'd47;
            32'h00000CC0: data = 32'd48;
            32'h00000CC4: data = 32'd49;
            32'h00000CC8: data = 32'd50;
            32'h00000CCC: data = 32'd51;
            32'h00000CD0: data = 32'd52;
            32'h00000CD4: data = 32'd53;
            32'h00000CD8: data = 32'd54;
            32'h00000CDC: data = 32'd55;
            32'h00000CE0: data = 32'd56;
            32'h00000CE4: data = 32'd57;
            32'h00000CE8: data = 32'd58;
            32'h00000CEC: data = 32'd59;
            32'h00000CF0: data = 32'd60;
            32'h00000CF4: data = 32'd61;
            32'h00000CF8: data = 32'd62;
            32'h00000CFC: data = 32'd63;
            32'h00000D00: data = 32'd64;
            32'h00000D04: data = 32'd65;
            32'h00000D08: data = 32'd66;
            32'h00000D0C: data = 32'd67;
            32'h00000D10: data = 32'd68;
            32'h00000D14: data = 32'd69;
            32'h00000D18: data = 32'd70;
            32'h00000D1C: data = 32'd71;
            32'h00000D20: data = 32'd72;
            32'h00000D24: data = 32'd73;
            32'h00000D28: data = 32'd74;
            32'h00000D2C: data = 32'd75;
            32'h00000D30: data = 32'd76;
            32'h00000D34: data = 32'd77;
            32'h00000D38: data = 32'd78;
            32'h00000D3C: data = 32'd79;
            32'h00000D40: data = 32'd80;
            32'h00000D44: data = 32'd81;
            32'h00000D48: data = 32'd82;
            32'h00000D4C: data = 32'd83;
            32'h00000D50: data = 32'd84;
            32'h00000D54: data = 32'd85;
            32'h00000D58: data = 32'd86;
            32'h00000D5C: data = 32'd87;
            32'h00000D60: data = 32'd88;
            32'h00000D64: data = 32'd89;
            32'h00000D68: data = 32'd90;
            32'h00000D6C: data = 32'd91;
            32'h00000D70: data = 32'd92;
            32'h00000D74: data = 32'd93;
            32'h00000D78: data = 32'd94;
            32'h00000D7C: data = 32'd95;
            32'h00000D80: data = 32'd96;
            32'h00000D84: data = 32'd97;
            32'h00000D88: data = 32'd98;
            32'h00000D8C: data = 32'd99;
            32'h00000D90: data = 32'd100;
            32'h00000D94: data = 32'd101;
            32'h00000D98: data = 32'd102;
            32'h00000D9C: data = 32'd103;
            32'h00000DA0: data = 32'd104;
            32'h00000DA4: data = 32'd105;
            32'h00000DA8: data = 32'd106;
            32'h00000DAC: data = 32'd107;
            32'h00000DB0: data = 32'd108;
            32'h00000DB4: data = 32'd109;
            32'h00000DB8: data = 32'd110;
            32'h00000DBC: data = 32'd111;
            32'h00000DC0: data = 32'd112;
            32'h00000DC4: data = 32'd113;
            32'h00000DC8: data = 32'd114;
            32'h00000DCC: data = 32'd115;
            32'h00000DD0: data = 32'd116;
            32'h00000DD4: data = 32'd117;
            32'h00000DD8: data = 32'd118;
            32'h00000DDC: data = 32'd119;
            32'h00000DE0: data = 32'd120;
            32'h00000DE4: data = 32'd121;
            32'h00000DE8: data = 32'd122;
            32'h00000DEC: data = 32'd123;
            32'h00000DF0: data = 32'd124;
            32'h00000DF4: data = 32'd125;
            32'h00000DF8: data = 32'd126;
            32'h00000DFC: data = 32'd127;
            32'h00000E00: data = 32'd128;
            32'h00000E04: data = 32'd129;
            32'h00000E08: data = 32'd130;
            32'h00000E0C: data = 32'd131;
            32'h00000E10: data = 32'd132;
            32'h00000E14: data = 32'd133;
            32'h00000E18: data = 32'd134;
            32'h00000E1C: data = 32'd135;
            32'h00000E20: data = 32'd136;
            32'h00000E24: data = 32'd137;
            32'h00000E28: data = 32'd138;
            32'h00000E2C: data = 32'd139;
            32'h00000E30: data = 32'd140;
            32'h00000E34: data = 32'd141;
            32'h00000E38: data = 32'd142;
            32'h00000E3C: data = 32'd143;
            32'h00000E40: data = 32'd144;
            32'h00000E44: data = 32'd145;
            32'h00000E48: data = 32'd146;
            32'h00000E4C: data = 32'd147;
            32'h00000E50: data = 32'd148;
            32'h00000E54: data = 32'd149;
            32'h00000E58: data = 32'd150;
            32'h00000E5C: data = 32'd151;
            32'h00000E60: data = 32'd152;
            32'h00000E64: data = 32'd153;
            32'h00000E68: data = 32'd154;
            32'h00000E6C: data = 32'd155;
            32'h00000E70: data = 32'd156;
            32'h00000E74: data = 32'd157;
            32'h00000E78: data = 32'd158;
            32'h00000E7C: data = 32'd159;
            32'h00000E80: data = 32'd160;
            32'h00000E84: data = 32'd161;
            32'h00000E88: data = 32'd162;
            32'h00000E8C: data = 32'd163;
            32'h00000E90: data = 32'd164;
            32'h00000E94: data = 32'd165;
            32'h00000E98: data = 32'd166;
            32'h00000E9C: data = 32'd167;
            32'h00000EA0: data = 32'd168;
            32'h00000EA4: data = 32'd169;
            32'h00000EA8: data = 32'd170;
            32'h00000EAC: data = 32'd171;
            32'h00000EB0: data = 32'd172;
            32'h00000EB4: data = 32'd173;
            32'h00000EB8: data = 32'd174;
            32'h00000EBC: data = 32'd175;
            32'h00000EC0: data = 32'd176;
            32'h00000EC4: data = 32'd177;
            32'h00000EC8: data = 32'd178;
            32'h00000ECC: data = 32'd179;
            32'h00000ED0: data = 32'd180;
            32'h00000ED4: data = 32'd181;
            32'h00000ED8: data = 32'd182;
            32'h00000EDC: data = 32'd183;
            32'h00000EE0: data = 32'd184;
            32'h00000EE4: data = 32'd185;
            32'h00000EE8: data = 32'd186;
            32'h00000EEC: data = 32'd187;
            32'h00000EF0: data = 32'd188;
            32'h00000EF4: data = 32'd189;
            32'h00000EF8: data = 32'd190;
            32'h00000EFC: data = 32'd191;
            32'h00000F00: data = 32'd192;
            32'h00000F04: data = 32'd193;
            32'h00000F08: data = 32'd194;
            32'h00000F0C: data = 32'd195;
            32'h00000F10: data = 32'd196;
            32'h00000F14: data = 32'd197;
            32'h00000F18: data = 32'd198;
            32'h00000F1C: data = 32'd199;
            32'h00000F20: data = 32'd200;
            32'h00000F24: data = 32'd201;
            32'h00000F28: data = 32'd202;
            32'h00000F2C: data = 32'd203;
            32'h00000F30: data = 32'd204;
            32'h00000F34: data = 32'd205;
            32'h00000F38: data = 32'd206;
            32'h00000F3C: data = 32'd207;
            32'h00000F40: data = 32'd208;
            32'h00000F44: data = 32'd209;
            32'h00000F48: data = 32'd210;
            32'h00000F4C: data = 32'd211;
            32'h00000F50: data = 32'd212;
            32'h00000F54: data = 32'd213;
            32'h00000F58: data = 32'd214;
            32'h00000F5C: data = 32'd215;
            32'h00000F60: data = 32'd216;
            32'h00000F64: data = 32'd217;
            32'h00000F68: data = 32'd218;
            32'h00000F6C: data = 32'd219;
            32'h00000F70: data = 32'd220;
            32'h00000F74: data = 32'd221;
            32'h00000F78: data = 32'd222;
            32'h00000F7C: data = 32'd223;
            32'h00000F80: data = 32'd224;
            32'h00000F84: data = 32'd225;
            32'h00000F88: data = 32'd226;
            32'h00000F8C: data = 32'd227;
            32'h00000F90: data = 32'd228;
            32'h00000F94: data = 32'd229;
            32'h00000F98: data = 32'd230;
            32'h00000F9C: data = 32'd231;
            32'h00000FA0: data = 32'd232;
            32'h00000FA4: data = 32'd233;
            32'h00000FA8: data = 32'd234;
            32'h00000FAC: data = 32'd235;
            32'h00000FB0: data = 32'd236;
            32'h00000FB4: data = 32'd237;
            32'h00000FB8: data = 32'd238;
            32'h00000FBC: data = 32'd239;
            32'h00000FC0: data = 32'd240;
            32'h00000FC4: data = 32'd241;
            32'h00000FC8: data = 32'd242;
            32'h00000FCC: data = 32'd243;
            32'h00000FD0: data = 32'd244;
            32'h00000FD4: data = 32'd245;
            32'h00000FD8: data = 32'd246;
            32'h00000FDC: data = 32'd247;
            32'h00000FE0: data = 32'd248;
            32'h00000FE4: data = 32'd249;
            32'h00000FE8: data = 32'd250;
            32'h00000FEC: data = 32'd251;
            32'h00000FF0: data = 32'd252;
            32'h00000FF4: data = 32'd253;
            32'h00000FF8: data = 32'd254;
            32'h00000FFC: data = 32'd255;
            32'h00001000: data = 32'd0;
            32'h00001004: data = 32'd1;
            32'h00001008: data = 32'd2;
            32'h0000100C: data = 32'd3;
            32'h00001010: data = 32'd4;
            32'h00001014: data = 32'd5;
            32'h00001018: data = 32'd6;
            32'h0000101C: data = 32'd7;
            32'h00001020: data = 32'd8;
            32'h00001024: data = 32'd9;
            32'h00001028: data = 32'd10;
            32'h0000102C: data = 32'd11;
            32'h00001030: data = 32'd12;
            32'h00001034: data = 32'd13;
            32'h00001038: data = 32'd14;
            32'h0000103C: data = 32'd15;
            32'h00001040: data = 32'd16;
            32'h00001044: data = 32'd17;
            32'h00001048: data = 32'd18;
            32'h0000104C: data = 32'd19;
            32'h00001050: data = 32'd20;
            32'h00001054: data = 32'd21;
            32'h00001058: data = 32'd22;
            32'h0000105C: data = 32'd23;
            32'h00001060: data = 32'd24;
            32'h00001064: data = 32'd25;
            32'h00001068: data = 32'd26;
            32'h0000106C: data = 32'd27;
            32'h00001070: data = 32'd28;
            32'h00001074: data = 32'd29;
            32'h00001078: data = 32'd30;
            32'h0000107C: data = 32'd31;
            32'h00001080: data = 32'd32;
            32'h00001084: data = 32'd33;
            32'h00001088: data = 32'd34;
            32'h0000108C: data = 32'd35;
            32'h00001090: data = 32'd36;
            32'h00001094: data = 32'd37;
            32'h00001098: data = 32'd38;
            32'h0000109C: data = 32'd39;
            32'h000010A0: data = 32'd40;
            32'h000010A4: data = 32'd41;
            32'h000010A8: data = 32'd42;
            32'h000010AC: data = 32'd43;
            32'h000010B0: data = 32'd44;
            32'h000010B4: data = 32'd45;
            32'h000010B8: data = 32'd46;
            32'h000010BC: data = 32'd47;
            32'h000010C0: data = 32'd48;
            32'h000010C4: data = 32'd49;
            32'h000010C8: data = 32'd50;
            32'h000010CC: data = 32'd51;
            32'h000010D0: data = 32'd52;
            32'h000010D4: data = 32'd53;
            32'h000010D8: data = 32'd54;
            32'h000010DC: data = 32'd55;
            32'h000010E0: data = 32'd56;
            32'h000010E4: data = 32'd57;
            32'h000010E8: data = 32'd58;
            32'h000010EC: data = 32'd59;
            32'h000010F0: data = 32'd60;
            32'h000010F4: data = 32'd61;
            32'h000010F8: data = 32'd62;
            32'h000010FC: data = 32'd63;
            32'h00001100: data = 32'd64;
            32'h00001104: data = 32'd65;
            32'h00001108: data = 32'd66;
            32'h0000110C: data = 32'd67;
            32'h00001110: data = 32'd68;
            32'h00001114: data = 32'd69;
            32'h00001118: data = 32'd70;
            32'h0000111C: data = 32'd71;
            32'h00001120: data = 32'd72;
            32'h00001124: data = 32'd73;
            32'h00001128: data = 32'd74;
            32'h0000112C: data = 32'd75;
            32'h00001130: data = 32'd76;
            32'h00001134: data = 32'd77;
            32'h00001138: data = 32'd78;
            32'h0000113C: data = 32'd79;
            32'h00001140: data = 32'd80;
            32'h00001144: data = 32'd81;
            32'h00001148: data = 32'd82;
            32'h0000114C: data = 32'd83;
            32'h00001150: data = 32'd84;
            32'h00001154: data = 32'd85;
            32'h00001158: data = 32'd86;
            32'h0000115C: data = 32'd87;
            32'h00001160: data = 32'd88;
            32'h00001164: data = 32'd89;
            32'h00001168: data = 32'd90;
            32'h0000116C: data = 32'd91;
            32'h00001170: data = 32'd92;
            32'h00001174: data = 32'd93;
            32'h00001178: data = 32'd94;
            32'h0000117C: data = 32'd95;
            32'h00001180: data = 32'd96;
            32'h00001184: data = 32'd97;
            32'h00001188: data = 32'd98;
            32'h0000118C: data = 32'd99;
            32'h00001190: data = 32'd100;
            32'h00001194: data = 32'd101;
            32'h00001198: data = 32'd102;
            32'h0000119C: data = 32'd103;
            32'h000011A0: data = 32'd104;
            32'h000011A4: data = 32'd105;
            32'h000011A8: data = 32'd106;
            32'h000011AC: data = 32'd107;
            32'h000011B0: data = 32'd108;
            32'h000011B4: data = 32'd109;
            32'h000011B8: data = 32'd110;
            32'h000011BC: data = 32'd111;
            32'h000011C0: data = 32'd112;
            32'h000011C4: data = 32'd113;
            32'h000011C8: data = 32'd114;
            32'h000011CC: data = 32'd115;
            32'h000011D0: data = 32'd116;
            32'h000011D4: data = 32'd117;
            32'h000011D8: data = 32'd118;
            32'h000011DC: data = 32'd119;
            32'h000011E0: data = 32'd120;
            32'h000011E4: data = 32'd121;
            32'h000011E8: data = 32'd122;
            32'h000011EC: data = 32'd123;
            32'h000011F0: data = 32'd124;
            32'h000011F4: data = 32'd125;
            32'h000011F8: data = 32'd126;
            32'h000011FC: data = 32'd127;
            32'h00001200: data = 32'd128;
            32'h00001204: data = 32'd129;
            32'h00001208: data = 32'd130;
            32'h0000120C: data = 32'd131;
            32'h00001210: data = 32'd132;
            32'h00001214: data = 32'd133;
            32'h00001218: data = 32'd134;
            32'h0000121C: data = 32'd135;
            32'h00001220: data = 32'd136;
            32'h00001224: data = 32'd137;
            32'h00001228: data = 32'd138;
            32'h0000122C: data = 32'd139;
            32'h00001230: data = 32'd140;
            32'h00001234: data = 32'd141;
            32'h00001238: data = 32'd142;
            32'h0000123C: data = 32'd143;
            32'h00001240: data = 32'd144;
            32'h00001244: data = 32'd145;
            32'h00001248: data = 32'd146;
            32'h0000124C: data = 32'd147;
            32'h00001250: data = 32'd148;
            32'h00001254: data = 32'd149;
            32'h00001258: data = 32'd150;
            32'h0000125C: data = 32'd151;
            32'h00001260: data = 32'd152;
            32'h00001264: data = 32'd153;
            32'h00001268: data = 32'd154;
            32'h0000126C: data = 32'd155;
            32'h00001270: data = 32'd156;
            32'h00001274: data = 32'd157;
            32'h00001278: data = 32'd158;
            32'h0000127C: data = 32'd159;
            32'h00001280: data = 32'd160;
            32'h00001284: data = 32'd161;
            32'h00001288: data = 32'd162;
            32'h0000128C: data = 32'd163;
            32'h00001290: data = 32'd164;
            32'h00001294: data = 32'd165;
            32'h00001298: data = 32'd166;
            32'h0000129C: data = 32'd167;
            32'h000012A0: data = 32'd168;
            32'h000012A4: data = 32'd169;
            32'h000012A8: data = 32'd170;
            32'h000012AC: data = 32'd171;
            32'h000012B0: data = 32'd172;
            32'h000012B4: data = 32'd173;
            32'h000012B8: data = 32'd174;
            32'h000012BC: data = 32'd175;
            32'h000012C0: data = 32'd176;
            32'h000012C4: data = 32'd177;
            32'h000012C8: data = 32'd178;
            32'h000012CC: data = 32'd179;
            32'h000012D0: data = 32'd180;
            32'h000012D4: data = 32'd181;
            32'h000012D8: data = 32'd182;
            32'h000012DC: data = 32'd183;
            32'h000012E0: data = 32'd184;
            32'h000012E4: data = 32'd185;
            32'h000012E8: data = 32'd186;
            32'h000012EC: data = 32'd187;
            32'h000012F0: data = 32'd188;
            32'h000012F4: data = 32'd189;
            32'h000012F8: data = 32'd190;
            32'h000012FC: data = 32'd191;
            32'h00001300: data = 32'd192;
            32'h00001304: data = 32'd193;
            32'h00001308: data = 32'd194;
            32'h0000130C: data = 32'd195;
            32'h00001310: data = 32'd196;
            32'h00001314: data = 32'd197;
            32'h00001318: data = 32'd198;
            32'h0000131C: data = 32'd199;
            32'h00001320: data = 32'd200;
            32'h00001324: data = 32'd201;
            32'h00001328: data = 32'd202;
            32'h0000132C: data = 32'd203;
            32'h00001330: data = 32'd204;
            32'h00001334: data = 32'd205;
            32'h00001338: data = 32'd206;
            32'h0000133C: data = 32'd207;
            32'h00001340: data = 32'd208;
            32'h00001344: data = 32'd209;
            32'h00001348: data = 32'd210;
            32'h0000134C: data = 32'd211;
            32'h00001350: data = 32'd212;
            32'h00001354: data = 32'd213;
            32'h00001358: data = 32'd214;
            32'h0000135C: data = 32'd215;
            32'h00001360: data = 32'd216;
            32'h00001364: data = 32'd217;
            32'h00001368: data = 32'd218;
            32'h0000136C: data = 32'd219;
            32'h00001370: data = 32'd220;
            32'h00001374: data = 32'd221;
            32'h00001378: data = 32'd222;
            32'h0000137C: data = 32'd223;
            32'h00001380: data = 32'd224;
            32'h00001384: data = 32'd225;
            32'h00001388: data = 32'd226;
            32'h0000138C: data = 32'd227;
            32'h00001390: data = 32'd228;
            32'h00001394: data = 32'd229;
            32'h00001398: data = 32'd230;
            32'h0000139C: data = 32'd231;
            32'h000013A0: data = 32'd232;
            32'h000013A4: data = 32'd233;
            32'h000013A8: data = 32'd234;
            32'h000013AC: data = 32'd235;
            32'h000013B0: data = 32'd236;
            32'h000013B4: data = 32'd237;
            32'h000013B8: data = 32'd238;
            32'h000013BC: data = 32'd239;
            32'h000013C0: data = 32'd240;
            32'h000013C4: data = 32'd241;
            32'h000013C8: data = 32'd242;
            32'h000013CC: data = 32'd243;
            32'h000013D0: data = 32'd244;
            32'h000013D4: data = 32'd245;
            32'h000013D8: data = 32'd246;
            32'h000013DC: data = 32'd247;
            32'h000013E0: data = 32'd248;
            32'h000013E4: data = 32'd249;
            32'h000013E8: data = 32'd250;
            32'h000013EC: data = 32'd251;
            32'h000013F0: data = 32'd252;
            32'h000013F4: data = 32'd253;
            32'h000013F8: data = 32'd254;
            32'h000013FC: data = 32'd255;
            32'h00001400: data = 32'd0;
            32'h00001404: data = 32'd1;
            32'h00001408: data = 32'd2;
            32'h0000140C: data = 32'd3;
            32'h00001410: data = 32'd4;
            32'h00001414: data = 32'd5;
            32'h00001418: data = 32'd6;
            32'h0000141C: data = 32'd7;
            32'h00001420: data = 32'd8;
            32'h00001424: data = 32'd9;
            32'h00001428: data = 32'd10;
            32'h0000142C: data = 32'd11;
            32'h00001430: data = 32'd12;
            32'h00001434: data = 32'd13;
            32'h00001438: data = 32'd14;
            32'h0000143C: data = 32'd15;
            32'h00001440: data = 32'd16;
            32'h00001444: data = 32'd17;
            32'h00001448: data = 32'd18;
            32'h0000144C: data = 32'd19;
            32'h00001450: data = 32'd20;
            32'h00001454: data = 32'd21;
            32'h00001458: data = 32'd22;
            32'h0000145C: data = 32'd23;
            32'h00001460: data = 32'd24;
            32'h00001464: data = 32'd25;
            32'h00001468: data = 32'd26;
            32'h0000146C: data = 32'd27;
            32'h00001470: data = 32'd28;
            32'h00001474: data = 32'd29;
            32'h00001478: data = 32'd30;
            32'h0000147C: data = 32'd31;
            32'h00001480: data = 32'd32;
            32'h00001484: data = 32'd33;
            32'h00001488: data = 32'd34;
            32'h0000148C: data = 32'd35;
            32'h00001490: data = 32'd36;
            32'h00001494: data = 32'd37;
            32'h00001498: data = 32'd38;
            32'h0000149C: data = 32'd39;
            32'h000014A0: data = 32'd40;
            32'h000014A4: data = 32'd41;
            32'h000014A8: data = 32'd42;
            32'h000014AC: data = 32'd43;
            32'h000014B0: data = 32'd44;
            32'h000014B4: data = 32'd45;
            32'h000014B8: data = 32'd46;
            32'h000014BC: data = 32'd47;
            32'h000014C0: data = 32'd48;
            32'h000014C4: data = 32'd49;
            32'h000014C8: data = 32'd50;
            32'h000014CC: data = 32'd51;
            32'h000014D0: data = 32'd52;
            32'h000014D4: data = 32'd53;
            32'h000014D8: data = 32'd54;
            32'h000014DC: data = 32'd55;
            32'h000014E0: data = 32'd56;
            32'h000014E4: data = 32'd57;
            32'h000014E8: data = 32'd58;
            32'h000014EC: data = 32'd59;
            32'h000014F0: data = 32'd60;
            32'h000014F4: data = 32'd61;
            32'h000014F8: data = 32'd62;
            32'h000014FC: data = 32'd63;
            32'h00001500: data = 32'd64;
            32'h00001504: data = 32'd65;
            32'h00001508: data = 32'd66;
            32'h0000150C: data = 32'd67;
            32'h00001510: data = 32'd68;
            32'h00001514: data = 32'd69;
            32'h00001518: data = 32'd70;
            32'h0000151C: data = 32'd71;
            32'h00001520: data = 32'd72;
            32'h00001524: data = 32'd73;
            32'h00001528: data = 32'd74;
            32'h0000152C: data = 32'd75;
            32'h00001530: data = 32'd76;
            32'h00001534: data = 32'd77;
            32'h00001538: data = 32'd78;
            32'h0000153C: data = 32'd79;
            32'h00001540: data = 32'd80;
            32'h00001544: data = 32'd81;
            32'h00001548: data = 32'd82;
            32'h0000154C: data = 32'd83;
            32'h00001550: data = 32'd84;
            32'h00001554: data = 32'd85;
            32'h00001558: data = 32'd86;
            32'h0000155C: data = 32'd87;
            32'h00001560: data = 32'd88;
            32'h00001564: data = 32'd89;
            32'h00001568: data = 32'd90;
            32'h0000156C: data = 32'd91;
            32'h00001570: data = 32'd92;
            32'h00001574: data = 32'd93;
            32'h00001578: data = 32'd94;
            32'h0000157C: data = 32'd95;
            32'h00001580: data = 32'd96;
            32'h00001584: data = 32'd97;
            32'h00001588: data = 32'd98;
            32'h0000158C: data = 32'd99;
            32'h00001590: data = 32'd100;
            32'h00001594: data = 32'd101;
            32'h00001598: data = 32'd102;
            32'h0000159C: data = 32'd103;
            32'h000015A0: data = 32'd104;
            32'h000015A4: data = 32'd105;
            32'h000015A8: data = 32'd106;
            32'h000015AC: data = 32'd107;
            32'h000015B0: data = 32'd108;
            32'h000015B4: data = 32'd109;
            32'h000015B8: data = 32'd110;
            32'h000015BC: data = 32'd111;
            32'h000015C0: data = 32'd112;
            32'h000015C4: data = 32'd113;
            32'h000015C8: data = 32'd114;
            32'h000015CC: data = 32'd115;
            32'h000015D0: data = 32'd116;
            32'h000015D4: data = 32'd117;
            32'h000015D8: data = 32'd118;
            32'h000015DC: data = 32'd119;
            32'h000015E0: data = 32'd120;
            32'h000015E4: data = 32'd121;
            32'h000015E8: data = 32'd122;
            32'h000015EC: data = 32'd123;
            32'h000015F0: data = 32'd124;
            32'h000015F4: data = 32'd125;
            32'h000015F8: data = 32'd126;
            32'h000015FC: data = 32'd127;
            32'h00001600: data = 32'd128;
            32'h00001604: data = 32'd129;
            32'h00001608: data = 32'd130;
            32'h0000160C: data = 32'd131;
            32'h00001610: data = 32'd132;
            32'h00001614: data = 32'd133;
            32'h00001618: data = 32'd134;
            32'h0000161C: data = 32'd135;
            32'h00001620: data = 32'd136;
            32'h00001624: data = 32'd137;
            32'h00001628: data = 32'd138;
            32'h0000162C: data = 32'd139;
            32'h00001630: data = 32'd140;
            32'h00001634: data = 32'd141;
            32'h00001638: data = 32'd142;
            32'h0000163C: data = 32'd143;
            32'h00001640: data = 32'd144;
            32'h00001644: data = 32'd145;
            32'h00001648: data = 32'd146;
            32'h0000164C: data = 32'd147;
            32'h00001650: data = 32'd148;
            32'h00001654: data = 32'd149;
            32'h00001658: data = 32'd150;
            32'h0000165C: data = 32'd151;
            32'h00001660: data = 32'd152;
            32'h00001664: data = 32'd153;
            32'h00001668: data = 32'd154;
            32'h0000166C: data = 32'd155;
            32'h00001670: data = 32'd156;
            32'h00001674: data = 32'd157;
            32'h00001678: data = 32'd158;
            32'h0000167C: data = 32'd159;
            32'h00001680: data = 32'd160;
            32'h00001684: data = 32'd161;
            32'h00001688: data = 32'd162;
            32'h0000168C: data = 32'd163;
            32'h00001690: data = 32'd164;
            32'h00001694: data = 32'd165;
            32'h00001698: data = 32'd166;
            32'h0000169C: data = 32'd167;
            32'h000016A0: data = 32'd168;
            32'h000016A4: data = 32'd169;
            32'h000016A8: data = 32'd170;
            32'h000016AC: data = 32'd171;
            32'h000016B0: data = 32'd172;
            32'h000016B4: data = 32'd173;
            32'h000016B8: data = 32'd174;
            32'h000016BC: data = 32'd175;
            32'h000016C0: data = 32'd176;
            32'h000016C4: data = 32'd177;
            32'h000016C8: data = 32'd178;
            32'h000016CC: data = 32'd179;
            32'h000016D0: data = 32'd180;
            32'h000016D4: data = 32'd181;
            32'h000016D8: data = 32'd182;
            32'h000016DC: data = 32'd183;
            32'h000016E0: data = 32'd184;
            32'h000016E4: data = 32'd185;
            32'h000016E8: data = 32'd186;
            32'h000016EC: data = 32'd187;
            32'h000016F0: data = 32'd188;
            32'h000016F4: data = 32'd189;
            32'h000016F8: data = 32'd190;
            32'h000016FC: data = 32'd191;
            32'h00001700: data = 32'd192;
            32'h00001704: data = 32'd193;
            32'h00001708: data = 32'd194;
            32'h0000170C: data = 32'd195;
            32'h00001710: data = 32'd196;
            32'h00001714: data = 32'd197;
            32'h00001718: data = 32'd198;
            32'h0000171C: data = 32'd199;
            32'h00001720: data = 32'd200;
            32'h00001724: data = 32'd201;
            32'h00001728: data = 32'd202;
            32'h0000172C: data = 32'd203;
            32'h00001730: data = 32'd204;
            32'h00001734: data = 32'd205;
            32'h00001738: data = 32'd206;
            32'h0000173C: data = 32'd207;
            32'h00001740: data = 32'd208;
            32'h00001744: data = 32'd209;
            32'h00001748: data = 32'd210;
            32'h0000174C: data = 32'd211;
            32'h00001750: data = 32'd212;
            32'h00001754: data = 32'd213;
            32'h00001758: data = 32'd214;
            32'h0000175C: data = 32'd215;
            32'h00001760: data = 32'd216;
            32'h00001764: data = 32'd217;
            32'h00001768: data = 32'd218;
            32'h0000176C: data = 32'd219;
            32'h00001770: data = 32'd220;
            32'h00001774: data = 32'd221;
            32'h00001778: data = 32'd222;
            32'h0000177C: data = 32'd223;
            32'h00001780: data = 32'd224;
            32'h00001784: data = 32'd225;
            32'h00001788: data = 32'd226;
            32'h0000178C: data = 32'd227;
            32'h00001790: data = 32'd228;
            32'h00001794: data = 32'd229;
            32'h00001798: data = 32'd230;
            32'h0000179C: data = 32'd231;
            32'h000017A0: data = 32'd232;
            32'h000017A4: data = 32'd233;
            32'h000017A8: data = 32'd234;
            32'h000017AC: data = 32'd235;
            32'h000017B0: data = 32'd236;
            32'h000017B4: data = 32'd237;
            32'h000017B8: data = 32'd238;
            32'h000017BC: data = 32'd239;
            32'h000017C0: data = 32'd240;
            32'h000017C4: data = 32'd241;
            32'h000017C8: data = 32'd242;
            32'h000017CC: data = 32'd243;
            32'h000017D0: data = 32'd244;
            32'h000017D4: data = 32'd245;
            32'h000017D8: data = 32'd246;
            32'h000017DC: data = 32'd247;
            32'h000017E0: data = 32'd248;
            32'h000017E4: data = 32'd249;
            32'h000017E8: data = 32'd250;
            32'h000017EC: data = 32'd251;
            32'h000017F0: data = 32'd252;
            32'h000017F4: data = 32'd253;
            32'h000017F8: data = 32'd254;
            32'h000017FC: data = 32'd255;
            32'h00001800: data = 32'd0;
            32'h00001804: data = 32'd1;
            32'h00001808: data = 32'd2;
            32'h0000180C: data = 32'd3;
            32'h00001810: data = 32'd4;
            32'h00001814: data = 32'd5;
            32'h00001818: data = 32'd6;
            32'h0000181C: data = 32'd7;
            32'h00001820: data = 32'd8;
            32'h00001824: data = 32'd9;
            32'h00001828: data = 32'd10;
            32'h0000182C: data = 32'd11;
            32'h00001830: data = 32'd12;
            32'h00001834: data = 32'd13;
            32'h00001838: data = 32'd14;
            32'h0000183C: data = 32'd15;
            32'h00001840: data = 32'd16;
            32'h00001844: data = 32'd17;
            32'h00001848: data = 32'd18;
            32'h0000184C: data = 32'd19;
            32'h00001850: data = 32'd20;
            32'h00001854: data = 32'd21;
            32'h00001858: data = 32'd22;
            32'h0000185C: data = 32'd23;
            32'h00001860: data = 32'd24;
            32'h00001864: data = 32'd25;
            32'h00001868: data = 32'd26;
            32'h0000186C: data = 32'd27;
            32'h00001870: data = 32'd28;
            32'h00001874: data = 32'd29;
            32'h00001878: data = 32'd30;
            32'h0000187C: data = 32'd31;
            32'h00001880: data = 32'd32;
            32'h00001884: data = 32'd33;
            32'h00001888: data = 32'd34;
            32'h0000188C: data = 32'd35;
            32'h00001890: data = 32'd36;
            32'h00001894: data = 32'd37;
            32'h00001898: data = 32'd38;
            32'h0000189C: data = 32'd39;
            32'h000018A0: data = 32'd40;
            32'h000018A4: data = 32'd41;
            32'h000018A8: data = 32'd42;
            32'h000018AC: data = 32'd43;
            32'h000018B0: data = 32'd44;
            32'h000018B4: data = 32'd45;
            32'h000018B8: data = 32'd46;
            32'h000018BC: data = 32'd47;
            32'h000018C0: data = 32'd48;
            32'h000018C4: data = 32'd49;
            32'h000018C8: data = 32'd50;
            32'h000018CC: data = 32'd51;
            32'h000018D0: data = 32'd52;
            32'h000018D4: data = 32'd53;
            32'h000018D8: data = 32'd54;
            32'h000018DC: data = 32'd55;
            32'h000018E0: data = 32'd56;
            32'h000018E4: data = 32'd57;
            32'h000018E8: data = 32'd58;
            32'h000018EC: data = 32'd59;
            32'h000018F0: data = 32'd60;
            32'h000018F4: data = 32'd61;
            32'h000018F8: data = 32'd62;
            32'h000018FC: data = 32'd63;
            32'h00001900: data = 32'd64;
            32'h00001904: data = 32'd65;
            32'h00001908: data = 32'd66;
            32'h0000190C: data = 32'd67;
            32'h00001910: data = 32'd68;
            32'h00001914: data = 32'd69;
            32'h00001918: data = 32'd70;
            32'h0000191C: data = 32'd71;
            32'h00001920: data = 32'd72;
            32'h00001924: data = 32'd73;
            32'h00001928: data = 32'd74;
            32'h0000192C: data = 32'd75;
            32'h00001930: data = 32'd76;
            32'h00001934: data = 32'd77;
            32'h00001938: data = 32'd78;
            32'h0000193C: data = 32'd79;
            32'h00001940: data = 32'd80;
            32'h00001944: data = 32'd81;
            32'h00001948: data = 32'd82;
            32'h0000194C: data = 32'd83;
            32'h00001950: data = 32'd84;
            32'h00001954: data = 32'd85;
            32'h00001958: data = 32'd86;
            32'h0000195C: data = 32'd87;
            32'h00001960: data = 32'd88;
            32'h00001964: data = 32'd89;
            32'h00001968: data = 32'd90;
            32'h0000196C: data = 32'd91;
            32'h00001970: data = 32'd92;
            32'h00001974: data = 32'd93;
            32'h00001978: data = 32'd94;
            32'h0000197C: data = 32'd95;
            32'h00001980: data = 32'd96;
            32'h00001984: data = 32'd97;
            32'h00001988: data = 32'd98;
            32'h0000198C: data = 32'd99;
            32'h00001990: data = 32'd100;
            32'h00001994: data = 32'd101;
            32'h00001998: data = 32'd102;
            32'h0000199C: data = 32'd103;
            32'h000019A0: data = 32'd104;
            32'h000019A4: data = 32'd105;
            32'h000019A8: data = 32'd106;
            32'h000019AC: data = 32'd107;
            32'h000019B0: data = 32'd108;
            32'h000019B4: data = 32'd109;
            32'h000019B8: data = 32'd110;
            32'h000019BC: data = 32'd111;
            32'h000019C0: data = 32'd112;
            32'h000019C4: data = 32'd113;
            32'h000019C8: data = 32'd114;
            32'h000019CC: data = 32'd115;
            32'h000019D0: data = 32'd116;
            32'h000019D4: data = 32'd117;
            32'h000019D8: data = 32'd118;
            32'h000019DC: data = 32'd119;
            32'h000019E0: data = 32'd120;
            32'h000019E4: data = 32'd121;
            32'h000019E8: data = 32'd122;
            32'h000019EC: data = 32'd123;
            32'h000019F0: data = 32'd124;
            32'h000019F4: data = 32'd125;
            32'h000019F8: data = 32'd126;
            32'h000019FC: data = 32'd127;
            32'h00001A00: data = 32'd128;
            32'h00001A04: data = 32'd129;
            32'h00001A08: data = 32'd130;
            32'h00001A0C: data = 32'd131;
            32'h00001A10: data = 32'd132;
            32'h00001A14: data = 32'd133;
            32'h00001A18: data = 32'd134;
            32'h00001A1C: data = 32'd135;
            32'h00001A20: data = 32'd136;
            32'h00001A24: data = 32'd137;
            32'h00001A28: data = 32'd138;
            32'h00001A2C: data = 32'd139;
            32'h00001A30: data = 32'd140;
            32'h00001A34: data = 32'd141;
            32'h00001A38: data = 32'd142;
            32'h00001A3C: data = 32'd143;
            32'h00001A40: data = 32'd144;
            32'h00001A44: data = 32'd145;
            32'h00001A48: data = 32'd146;
            32'h00001A4C: data = 32'd147;
            32'h00001A50: data = 32'd148;
            32'h00001A54: data = 32'd149;
            32'h00001A58: data = 32'd150;
            32'h00001A5C: data = 32'd151;
            32'h00001A60: data = 32'd152;
            32'h00001A64: data = 32'd153;
            32'h00001A68: data = 32'd154;
            32'h00001A6C: data = 32'd155;
            32'h00001A70: data = 32'd156;
            32'h00001A74: data = 32'd157;
            32'h00001A78: data = 32'd158;
            32'h00001A7C: data = 32'd159;
            32'h00001A80: data = 32'd160;
            32'h00001A84: data = 32'd161;
            32'h00001A88: data = 32'd162;
            32'h00001A8C: data = 32'd163;
            32'h00001A90: data = 32'd164;
            32'h00001A94: data = 32'd165;
            32'h00001A98: data = 32'd166;
            32'h00001A9C: data = 32'd167;
            32'h00001AA0: data = 32'd168;
            32'h00001AA4: data = 32'd169;
            32'h00001AA8: data = 32'd170;
            32'h00001AAC: data = 32'd171;
            32'h00001AB0: data = 32'd172;
            32'h00001AB4: data = 32'd173;
            32'h00001AB8: data = 32'd174;
            32'h00001ABC: data = 32'd175;
            32'h00001AC0: data = 32'd176;
            32'h00001AC4: data = 32'd177;
            32'h00001AC8: data = 32'd178;
            32'h00001ACC: data = 32'd179;
            32'h00001AD0: data = 32'd180;
            32'h00001AD4: data = 32'd181;
            32'h00001AD8: data = 32'd182;
            32'h00001ADC: data = 32'd183;
            32'h00001AE0: data = 32'd184;
            32'h00001AE4: data = 32'd185;
            32'h00001AE8: data = 32'd186;
            32'h00001AEC: data = 32'd187;
            32'h00001AF0: data = 32'd188;
            32'h00001AF4: data = 32'd189;
            32'h00001AF8: data = 32'd190;
            32'h00001AFC: data = 32'd191;
            32'h00001B00: data = 32'd192;
            32'h00001B04: data = 32'd193;
            32'h00001B08: data = 32'd194;
            32'h00001B0C: data = 32'd195;
            32'h00001B10: data = 32'd196;
            32'h00001B14: data = 32'd197;
            32'h00001B18: data = 32'd198;
            32'h00001B1C: data = 32'd199;
            32'h00001B20: data = 32'd200;
            32'h00001B24: data = 32'd201;
            32'h00001B28: data = 32'd202;
            32'h00001B2C: data = 32'd203;
            32'h00001B30: data = 32'd204;
            32'h00001B34: data = 32'd205;
            32'h00001B38: data = 32'd206;
            32'h00001B3C: data = 32'd207;
            32'h00001B40: data = 32'd208;
            32'h00001B44: data = 32'd209;
            32'h00001B48: data = 32'd210;
            32'h00001B4C: data = 32'd211;
            32'h00001B50: data = 32'd212;
            32'h00001B54: data = 32'd213;
            32'h00001B58: data = 32'd214;
            32'h00001B5C: data = 32'd215;
            32'h00001B60: data = 32'd216;
            32'h00001B64: data = 32'd217;
            32'h00001B68: data = 32'd218;
            32'h00001B6C: data = 32'd219;
            32'h00001B70: data = 32'd220;
            32'h00001B74: data = 32'd221;
            32'h00001B78: data = 32'd222;
            32'h00001B7C: data = 32'd223;
            32'h00001B80: data = 32'd224;
            32'h00001B84: data = 32'd225;
            32'h00001B88: data = 32'd226;
            32'h00001B8C: data = 32'd227;
            32'h00001B90: data = 32'd228;
            32'h00001B94: data = 32'd229;
            32'h00001B98: data = 32'd230;
            32'h00001B9C: data = 32'd231;
            32'h00001BA0: data = 32'd232;
            32'h00001BA4: data = 32'd233;
            32'h00001BA8: data = 32'd234;
            32'h00001BAC: data = 32'd235;
            32'h00001BB0: data = 32'd236;
            32'h00001BB4: data = 32'd237;
            32'h00001BB8: data = 32'd238;
            32'h00001BBC: data = 32'd239;
            32'h00001BC0: data = 32'd240;
            32'h00001BC4: data = 32'd241;
            32'h00001BC8: data = 32'd242;
            32'h00001BCC: data = 32'd243;
            32'h00001BD0: data = 32'd244;
            32'h00001BD4: data = 32'd245;
            32'h00001BD8: data = 32'd246;
            32'h00001BDC: data = 32'd247;
            32'h00001BE0: data = 32'd248;
            32'h00001BE4: data = 32'd249;
            32'h00001BE8: data = 32'd250;
            32'h00001BEC: data = 32'd251;
            32'h00001BF0: data = 32'd252;
            32'h00001BF4: data = 32'd253;
            32'h00001BF8: data = 32'd254;
            32'h00001BFC: data = 32'd255;
            32'h00001C00: data = 32'd0;
            32'h00001C04: data = 32'd1;
            32'h00001C08: data = 32'd2;
            32'h00001C0C: data = 32'd3;
            32'h00001C10: data = 32'd4;
            32'h00001C14: data = 32'd5;
            32'h00001C18: data = 32'd6;
            32'h00001C1C: data = 32'd7;
            32'h00001C20: data = 32'd8;
            32'h00001C24: data = 32'd9;
            32'h00001C28: data = 32'd10;
            32'h00001C2C: data = 32'd11;
            32'h00001C30: data = 32'd12;
            32'h00001C34: data = 32'd13;
            32'h00001C38: data = 32'd14;
            32'h00001C3C: data = 32'd15;
            32'h00001C40: data = 32'd16;
            32'h00001C44: data = 32'd17;
            32'h00001C48: data = 32'd18;
            32'h00001C4C: data = 32'd19;
            32'h00001C50: data = 32'd20;
            32'h00001C54: data = 32'd21;
            32'h00001C58: data = 32'd22;
            32'h00001C5C: data = 32'd23;
            32'h00001C60: data = 32'd24;
            32'h00001C64: data = 32'd25;
            32'h00001C68: data = 32'd26;
            32'h00001C6C: data = 32'd27;
            32'h00001C70: data = 32'd28;
            32'h00001C74: data = 32'd29;
            32'h00001C78: data = 32'd30;
            32'h00001C7C: data = 32'd31;
            32'h00001C80: data = 32'd32;
            32'h00001C84: data = 32'd33;
            32'h00001C88: data = 32'd34;
            32'h00001C8C: data = 32'd35;
            32'h00001C90: data = 32'd36;
            32'h00001C94: data = 32'd37;
            32'h00001C98: data = 32'd38;
            32'h00001C9C: data = 32'd39;
            32'h00001CA0: data = 32'd40;
            32'h00001CA4: data = 32'd41;
            32'h00001CA8: data = 32'd42;
            32'h00001CAC: data = 32'd43;
            32'h00001CB0: data = 32'd44;
            32'h00001CB4: data = 32'd45;
            32'h00001CB8: data = 32'd46;
            32'h00001CBC: data = 32'd47;
            32'h00001CC0: data = 32'd48;
            32'h00001CC4: data = 32'd49;
            32'h00001CC8: data = 32'd50;
            32'h00001CCC: data = 32'd51;
            32'h00001CD0: data = 32'd52;
            32'h00001CD4: data = 32'd53;
            32'h00001CD8: data = 32'd54;
            32'h00001CDC: data = 32'd55;
            32'h00001CE0: data = 32'd56;
            32'h00001CE4: data = 32'd57;
            32'h00001CE8: data = 32'd58;
            32'h00001CEC: data = 32'd59;
            32'h00001CF0: data = 32'd60;
            32'h00001CF4: data = 32'd61;
            32'h00001CF8: data = 32'd62;
            32'h00001CFC: data = 32'd63;
            32'h00001D00: data = 32'd64;
            32'h00001D04: data = 32'd65;
            32'h00001D08: data = 32'd66;
            32'h00001D0C: data = 32'd67;
            32'h00001D10: data = 32'd68;
            32'h00001D14: data = 32'd69;
            32'h00001D18: data = 32'd70;
            32'h00001D1C: data = 32'd71;
            32'h00001D20: data = 32'd72;
            32'h00001D24: data = 32'd73;
            32'h00001D28: data = 32'd74;
            32'h00001D2C: data = 32'd75;
            32'h00001D30: data = 32'd76;
            32'h00001D34: data = 32'd77;
            32'h00001D38: data = 32'd78;
            32'h00001D3C: data = 32'd79;
            32'h00001D40: data = 32'd80;
            32'h00001D44: data = 32'd81;
            32'h00001D48: data = 32'd82;
            32'h00001D4C: data = 32'd83;
            32'h00001D50: data = 32'd84;
            32'h00001D54: data = 32'd85;
            32'h00001D58: data = 32'd86;
            32'h00001D5C: data = 32'd87;
            32'h00001D60: data = 32'd88;
            32'h00001D64: data = 32'd89;
            32'h00001D68: data = 32'd90;
            32'h00001D6C: data = 32'd91;
            32'h00001D70: data = 32'd92;
            32'h00001D74: data = 32'd93;
            32'h00001D78: data = 32'd94;
            32'h00001D7C: data = 32'd95;
            32'h00001D80: data = 32'd96;
            32'h00001D84: data = 32'd97;
            32'h00001D88: data = 32'd98;
            32'h00001D8C: data = 32'd99;
            32'h00001D90: data = 32'd100;
            32'h00001D94: data = 32'd101;
            32'h00001D98: data = 32'd102;
            32'h00001D9C: data = 32'd103;
            32'h00001DA0: data = 32'd104;
            32'h00001DA4: data = 32'd105;
            32'h00001DA8: data = 32'd106;
            32'h00001DAC: data = 32'd107;
            32'h00001DB0: data = 32'd108;
            32'h00001DB4: data = 32'd109;
            32'h00001DB8: data = 32'd110;
            32'h00001DBC: data = 32'd111;
            32'h00001DC0: data = 32'd112;
            32'h00001DC4: data = 32'd113;
            32'h00001DC8: data = 32'd114;
            32'h00001DCC: data = 32'd115;
            32'h00001DD0: data = 32'd116;
            32'h00001DD4: data = 32'd117;
            32'h00001DD8: data = 32'd118;
            32'h00001DDC: data = 32'd119;
            32'h00001DE0: data = 32'd120;
            32'h00001DE4: data = 32'd121;
            32'h00001DE8: data = 32'd122;
            32'h00001DEC: data = 32'd123;
            32'h00001DF0: data = 32'd124;
            32'h00001DF4: data = 32'd125;
            32'h00001DF8: data = 32'd126;
            32'h00001DFC: data = 32'd127;
            32'h00001E00: data = 32'd128;
            32'h00001E04: data = 32'd129;
            32'h00001E08: data = 32'd130;
            32'h00001E0C: data = 32'd131;
            32'h00001E10: data = 32'd132;
            32'h00001E14: data = 32'd133;
            32'h00001E18: data = 32'd134;
            32'h00001E1C: data = 32'd135;
            32'h00001E20: data = 32'd136;
            32'h00001E24: data = 32'd137;
            32'h00001E28: data = 32'd138;
            32'h00001E2C: data = 32'd139;
            32'h00001E30: data = 32'd140;
            32'h00001E34: data = 32'd141;
            32'h00001E38: data = 32'd142;
            32'h00001E3C: data = 32'd143;
            32'h00001E40: data = 32'd144;
            32'h00001E44: data = 32'd145;
            32'h00001E48: data = 32'd146;
            32'h00001E4C: data = 32'd147;
            32'h00001E50: data = 32'd148;
            32'h00001E54: data = 32'd149;
            32'h00001E58: data = 32'd150;
            32'h00001E5C: data = 32'd151;
            32'h00001E60: data = 32'd152;
            32'h00001E64: data = 32'd153;
            32'h00001E68: data = 32'd154;
            32'h00001E6C: data = 32'd155;
            32'h00001E70: data = 32'd156;
            32'h00001E74: data = 32'd157;
            32'h00001E78: data = 32'd158;
            32'h00001E7C: data = 32'd159;
            32'h00001E80: data = 32'd160;
            32'h00001E84: data = 32'd161;
            32'h00001E88: data = 32'd162;
            32'h00001E8C: data = 32'd163;
            32'h00001E90: data = 32'd164;
            32'h00001E94: data = 32'd165;
            32'h00001E98: data = 32'd166;
            32'h00001E9C: data = 32'd167;
            32'h00001EA0: data = 32'd168;
            32'h00001EA4: data = 32'd169;
            32'h00001EA8: data = 32'd170;
            32'h00001EAC: data = 32'd171;
            32'h00001EB0: data = 32'd172;
            32'h00001EB4: data = 32'd173;
            32'h00001EB8: data = 32'd174;
            32'h00001EBC: data = 32'd175;
            32'h00001EC0: data = 32'd176;
            32'h00001EC4: data = 32'd177;
            32'h00001EC8: data = 32'd178;
            32'h00001ECC: data = 32'd179;
            32'h00001ED0: data = 32'd180;
            32'h00001ED4: data = 32'd181;
            32'h00001ED8: data = 32'd182;
            32'h00001EDC: data = 32'd183;
            32'h00001EE0: data = 32'd184;
            32'h00001EE4: data = 32'd185;
            32'h00001EE8: data = 32'd186;
            32'h00001EEC: data = 32'd187;
            32'h00001EF0: data = 32'd188;
            32'h00001EF4: data = 32'd189;
            32'h00001EF8: data = 32'd190;
            32'h00001EFC: data = 32'd191;
            32'h00001F00: data = 32'd192;
            32'h00001F04: data = 32'd193;
            32'h00001F08: data = 32'd194;
            32'h00001F0C: data = 32'd195;
            32'h00001F10: data = 32'd196;
            32'h00001F14: data = 32'd197;
            32'h00001F18: data = 32'd198;
            32'h00001F1C: data = 32'd199;
            32'h00001F20: data = 32'd200;
            32'h00001F24: data = 32'd201;
            32'h00001F28: data = 32'd202;
            32'h00001F2C: data = 32'd203;
            32'h00001F30: data = 32'd204;
            32'h00001F34: data = 32'd205;
            32'h00001F38: data = 32'd206;
            32'h00001F3C: data = 32'd207;
            default: data = 32'd0;
        endcase
    end

endmodule

