

module BRAM_sim_biiiig (
    input  logic [31:0] address,
    output logic [31:0]  data_send,
    input logic clk,
    input logic reset
);
    logic [31:0] data;
    
    always_ff @(posedge clk)
    if (reset)
    data_send <= 32'd0;
    else
    data_send <= data;



    always_comb begin
        case (address)
            32'hB0000000: data = 32'd0;
            32'hB0000004: data = 32'd1;
            32'hB0000008: data = 32'd2;
            32'hB000000C: data = 32'd3;
            32'hB0000010: data = 32'd4;
            32'hB0000014: data = 32'd5;
            32'hB0000018: data = 32'd6;
            32'hB000001C: data = 32'd7;
            32'hB0000020: data = 32'd8;
            32'hB0000024: data = 32'd9;
            32'hB0000028: data = 32'd10;
            32'hB000002C: data = 32'd11;
            32'hB0000030: data = 32'd12;
            32'hB0000034: data = 32'd13;
            32'hB0000038: data = 32'd14;
            32'hB000003C: data = 32'd15;
            32'hB0000040: data = 32'd16;
            32'hB0000044: data = 32'd17;
            32'hB0000048: data = 32'd18;
            32'hB000004C: data = 32'd19;
            32'hB0000050: data = 32'd20;
            32'hB0000054: data = 32'd21;
            32'hB0000058: data = 32'd22;
            32'hB000005C: data = 32'd23;
            32'hB0000060: data = 32'd24;
            32'hB0000064: data = 32'd25;
            32'hB0000068: data = 32'd26;
            32'hB000006C: data = 32'd27;
            32'hB0000070: data = 32'd28;
            32'hB0000074: data = 32'd29;
            32'hB0000078: data = 32'd30;
            32'hB000007C: data = 32'd31;
            32'hB0000080: data = 32'd32;
            32'hB0000084: data = 32'd33;
            32'hB0000088: data = 32'd34;
            32'hB000008C: data = 32'd35;
            32'hB0000090: data = 32'd36;
            32'hB0000094: data = 32'd37;
            32'hB0000098: data = 32'd38;
            32'hB000009C: data = 32'd39;
            32'hB00000A0: data = 32'd40;
            32'hB00000A4: data = 32'd41;
            32'hB00000A8: data = 32'd42;
            32'hB00000AC: data = 32'd43;
            32'hB00000B0: data = 32'd44;
            32'hB00000B4: data = 32'd45;
            32'hB00000B8: data = 32'd46;
            32'hB00000BC: data = 32'd47;
            32'hB00000C0: data = 32'd48;
            32'hB00000C4: data = 32'd49;
            32'hB00000C8: data = 32'd50;
            32'hB00000CC: data = 32'd51;
            32'hB00000D0: data = 32'd52;
            32'hB00000D4: data = 32'd53;
            32'hB00000D8: data = 32'd54;
            32'hB00000DC: data = 32'd55;
            32'hB00000E0: data = 32'd56;
            32'hB00000E4: data = 32'd57;
            32'hB00000E8: data = 32'd58;
            32'hB00000EC: data = 32'd59;
            32'hB00000F0: data = 32'd60;
            32'hB00000F4: data = 32'd61;
            32'hB00000F8: data = 32'd62;
            32'hB00000FC: data = 32'd63;
            32'hB0000100: data = 32'd64;
            32'hB0000104: data = 32'd65;
            32'hB0000108: data = 32'd66;
            32'hB000010C: data = 32'd67;
            32'hB0000110: data = 32'd68;
            32'hB0000114: data = 32'd69;
            32'hB0000118: data = 32'd70;
            32'hB000011C: data = 32'd71;
            32'hB0000120: data = 32'd72;
            32'hB0000124: data = 32'd73;
            32'hB0000128: data = 32'd74;
            32'hB000012C: data = 32'd75;
            32'hB0000130: data = 32'd76;
            32'hB0000134: data = 32'd77;
            32'hB0000138: data = 32'd78;
            32'hB000013C: data = 32'd79;
            32'hB0000140: data = 32'd80;
            32'hB0000144: data = 32'd81;
            32'hB0000148: data = 32'd82;
            32'hB000014C: data = 32'd83;
            32'hB0000150: data = 32'd84;
            32'hB0000154: data = 32'd85;
            32'hB0000158: data = 32'd86;
            32'hB000015C: data = 32'd87;
            32'hB0000160: data = 32'd88;
            32'hB0000164: data = 32'd89;
            32'hB0000168: data = 32'd90;
            32'hB000016C: data = 32'd91;
            32'hB0000170: data = 32'd92;
            32'hB0000174: data = 32'd93;
            32'hB0000178: data = 32'd94;
            32'hB000017C: data = 32'd95;
            32'hB0000180: data = 32'd96;
            32'hB0000184: data = 32'd97;
            32'hB0000188: data = 32'd98;
            32'hB000018C: data = 32'd99;
            32'hB0000190: data = 32'd100;
            32'hB0000194: data = 32'd101;
            32'hB0000198: data = 32'd102;
            32'hB000019C: data = 32'd103;
            32'hB00001A0: data = 32'd104;
            32'hB00001A4: data = 32'd105;
            32'hB00001A8: data = 32'd106;
            32'hB00001AC: data = 32'd107;
            32'hB00001B0: data = 32'd108;
            32'hB00001B4: data = 32'd109;
            32'hB00001B8: data = 32'd110;
            32'hB00001BC: data = 32'd111;
            32'hB00001C0: data = 32'd112;
            32'hB00001C4: data = 32'd113;
            32'hB00001C8: data = 32'd114;
            32'hB00001CC: data = 32'd115;
            32'hB00001D0: data = 32'd116;
            32'hB00001D4: data = 32'd117;
            32'hB00001D8: data = 32'd118;
            32'hB00001DC: data = 32'd119;
            32'hB00001E0: data = 32'd120;
            32'hB00001E4: data = 32'd121;
            32'hB00001E8: data = 32'd122;
            32'hB00001EC: data = 32'd123;
            32'hB00001F0: data = 32'd124;
            32'hB00001F4: data = 32'd125;
            32'hB00001F8: data = 32'd126;
            32'hB00001FC: data = 32'd127;
            32'hB0000200: data = 32'd128;
            32'hB0000204: data = 32'd129;
            32'hB0000208: data = 32'd130;
            32'hB000020C: data = 32'd131;
            32'hB0000210: data = 32'd132;
            32'hB0000214: data = 32'd133;
            32'hB0000218: data = 32'd134;
            32'hB000021C: data = 32'd135;
            32'hB0000220: data = 32'd136;
            32'hB0000224: data = 32'd137;
            32'hB0000228: data = 32'd138;
            32'hB000022C: data = 32'd139;
            32'hB0000230: data = 32'd140;
            32'hB0000234: data = 32'd141;
            32'hB0000238: data = 32'd142;
            32'hB000023C: data = 32'd143;
            32'hB0000240: data = 32'd144;
            32'hB0000244: data = 32'd145;
            32'hB0000248: data = 32'd146;
            32'hB000024C: data = 32'd147;
            32'hB0000250: data = 32'd148;
            32'hB0000254: data = 32'd149;
            32'hB0000258: data = 32'd150;
            32'hB000025C: data = 32'd151;
            32'hB0000260: data = 32'd152;
            32'hB0000264: data = 32'd153;
            32'hB0000268: data = 32'd154;
            32'hB000026C: data = 32'd155;
            32'hB0000270: data = 32'd156;
            32'hB0000274: data = 32'd157;
            32'hB0000278: data = 32'd158;
            32'hB000027C: data = 32'd159;
            32'hB0000280: data = 32'd160;
            32'hB0000284: data = 32'd161;
            32'hB0000288: data = 32'd162;
            32'hB000028C: data = 32'd163;
            32'hB0000290: data = 32'd164;
            32'hB0000294: data = 32'd165;
            32'hB0000298: data = 32'd166;
            32'hB000029C: data = 32'd167;
            32'hB00002A0: data = 32'd168;
            32'hB00002A4: data = 32'd169;
            32'hB00002A8: data = 32'd170;
            32'hB00002AC: data = 32'd171;
            32'hB00002B0: data = 32'd172;
            32'hB00002B4: data = 32'd173;
            32'hB00002B8: data = 32'd174;
            32'hB00002BC: data = 32'd175;
            32'hB00002C0: data = 32'd176;
            32'hB00002C4: data = 32'd177;
            32'hB00002C8: data = 32'd178;
            32'hB00002CC: data = 32'd179;
            32'hB00002D0: data = 32'd180;
            32'hB00002D4: data = 32'd181;
            32'hB00002D8: data = 32'd182;
            32'hB00002DC: data = 32'd183;
            32'hB00002E0: data = 32'd184;
            32'hB00002E4: data = 32'd185;
            32'hB00002E8: data = 32'd186;
            32'hB00002EC: data = 32'd187;
            32'hB00002F0: data = 32'd188;
            32'hB00002F4: data = 32'd189;
            32'hB00002F8: data = 32'd190;
            32'hB00002FC: data = 32'd191;
            32'hB0000300: data = 32'd192;
            32'hB0000304: data = 32'd193;
            32'hB0000308: data = 32'd194;
            32'hB000030C: data = 32'd195;
            32'hB0000310: data = 32'd196;
            32'hB0000314: data = 32'd197;
            32'hB0000318: data = 32'd198;
            32'hB000031C: data = 32'd199;
            32'hB0000320: data = 32'd200;
            32'hB0000324: data = 32'd201;
            32'hB0000328: data = 32'd202;
            32'hB000032C: data = 32'd203;
            32'hB0000330: data = 32'd204;
            32'hB0000334: data = 32'd205;
            32'hB0000338: data = 32'd206;
            32'hB000033C: data = 32'd207;
            32'hB0000340: data = 32'd208;
            32'hB0000344: data = 32'd209;
            32'hB0000348: data = 32'd210;
            32'hB000034C: data = 32'd211;
            32'hB0000350: data = 32'd212;
            32'hB0000354: data = 32'd213;
            32'hB0000358: data = 32'd214;
            32'hB000035C: data = 32'd215;
            32'hB0000360: data = 32'd216;
            32'hB0000364: data = 32'd217;
            32'hB0000368: data = 32'd218;
            32'hB000036C: data = 32'd219;
            32'hB0000370: data = 32'd220;
            32'hB0000374: data = 32'd221;
            32'hB0000378: data = 32'd222;
            32'hB000037C: data = 32'd223;
            32'hB0000380: data = 32'd224;
            32'hB0000384: data = 32'd225;
            32'hB0000388: data = 32'd226;
            32'hB000038C: data = 32'd227;
            32'hB0000390: data = 32'd228;
            32'hB0000394: data = 32'd229;
            32'hB0000398: data = 32'd230;
            32'hB000039C: data = 32'd231;
            32'hB00003A0: data = 32'd232;
            32'hB00003A4: data = 32'd233;
            32'hB00003A8: data = 32'd234;
            32'hB00003AC: data = 32'd235;
            32'hB00003B0: data = 32'd236;
            32'hB00003B4: data = 32'd237;
            32'hB00003B8: data = 32'd238;
            32'hB00003BC: data = 32'd239;
            32'hB00003C0: data = 32'd240;
            32'hB00003C4: data = 32'd241;
            32'hB00003C8: data = 32'd242;
            32'hB00003CC: data = 32'd243;
            32'hB00003D0: data = 32'd244;
            32'hB00003D4: data = 32'd245;
            32'hB00003D8: data = 32'd246;
            32'hB00003DC: data = 32'd247;
            32'hB00003E0: data = 32'd248;
            32'hB00003E4: data = 32'd249;
            32'hB00003E8: data = 32'd250;
            32'hB00003EC: data = 32'd251;
            32'hB00003F0: data = 32'd252;
            32'hB00003F4: data = 32'd253;
            32'hB00003F8: data = 32'd254;
            32'hB00003FC: data = 32'd255;
            32'hB0000400: data = 32'd0;
            32'hB0000404: data = 32'd1;
            32'hB0000408: data = 32'd2;
            32'hB000040C: data = 32'd3;
            32'hB0000410: data = 32'd4;
            32'hB0000414: data = 32'd5;
            32'hB0000418: data = 32'd6;
            32'hB000041C: data = 32'd7;
            32'hB0000420: data = 32'd8;
            32'hB0000424: data = 32'd9;
            32'hB0000428: data = 32'd10;
            32'hB000042C: data = 32'd11;
            32'hB0000430: data = 32'd12;
            32'hB0000434: data = 32'd13;
            32'hB0000438: data = 32'd14;
            32'hB000043C: data = 32'd15;
            32'hB0000440: data = 32'd16;
            32'hB0000444: data = 32'd17;
            32'hB0000448: data = 32'd18;
            32'hB000044C: data = 32'd19;
            32'hB0000450: data = 32'd20;
            32'hB0000454: data = 32'd21;
            32'hB0000458: data = 32'd22;
            32'hB000045C: data = 32'd23;
            32'hB0000460: data = 32'd24;
            32'hB0000464: data = 32'd25;
            32'hB0000468: data = 32'd26;
            32'hB000046C: data = 32'd27;
            32'hB0000470: data = 32'd28;
            32'hB0000474: data = 32'd29;
            32'hB0000478: data = 32'd30;
            32'hB000047C: data = 32'd31;
            32'hB0000480: data = 32'd32;
            32'hB0000484: data = 32'd33;
            32'hB0000488: data = 32'd34;
            32'hB000048C: data = 32'd35;
            32'hB0000490: data = 32'd36;
            32'hB0000494: data = 32'd37;
            32'hB0000498: data = 32'd38;
            32'hB000049C: data = 32'd39;
            32'hB00004A0: data = 32'd40;
            32'hB00004A4: data = 32'd41;
            32'hB00004A8: data = 32'd42;
            32'hB00004AC: data = 32'd43;
            32'hB00004B0: data = 32'd44;
            32'hB00004B4: data = 32'd45;
            32'hB00004B8: data = 32'd46;
            32'hB00004BC: data = 32'd47;
            32'hB00004C0: data = 32'd48;
            32'hB00004C4: data = 32'd49;
            32'hB00004C8: data = 32'd50;
            32'hB00004CC: data = 32'd51;
            32'hB00004D0: data = 32'd52;
            32'hB00004D4: data = 32'd53;
            32'hB00004D8: data = 32'd54;
            32'hB00004DC: data = 32'd55;
            32'hB00004E0: data = 32'd56;
            32'hB00004E4: data = 32'd57;
            32'hB00004E8: data = 32'd58;
            32'hB00004EC: data = 32'd59;
            32'hB00004F0: data = 32'd60;
            32'hB00004F4: data = 32'd61;
            32'hB00004F8: data = 32'd62;
            32'hB00004FC: data = 32'd63;
            32'hB0000500: data = 32'd64;
            32'hB0000504: data = 32'd65;
            32'hB0000508: data = 32'd66;
            32'hB000050C: data = 32'd67;
            32'hB0000510: data = 32'd68;
            32'hB0000514: data = 32'd69;
            32'hB0000518: data = 32'd70;
            32'hB000051C: data = 32'd71;
            32'hB0000520: data = 32'd72;
            32'hB0000524: data = 32'd73;
            32'hB0000528: data = 32'd74;
            32'hB000052C: data = 32'd75;
            32'hB0000530: data = 32'd76;
            32'hB0000534: data = 32'd77;
            32'hB0000538: data = 32'd78;
            32'hB000053C: data = 32'd79;
            32'hB0000540: data = 32'd80;
            32'hB0000544: data = 32'd81;
            32'hB0000548: data = 32'd82;
            32'hB000054C: data = 32'd83;
            32'hB0000550: data = 32'd84;
            32'hB0000554: data = 32'd85;
            32'hB0000558: data = 32'd86;
            32'hB000055C: data = 32'd87;
            32'hB0000560: data = 32'd88;
            32'hB0000564: data = 32'd89;
            32'hB0000568: data = 32'd90;
            32'hB000056C: data = 32'd91;
            32'hB0000570: data = 32'd92;
            32'hB0000574: data = 32'd93;
            32'hB0000578: data = 32'd94;
            32'hB000057C: data = 32'd95;
            32'hB0000580: data = 32'd96;
            32'hB0000584: data = 32'd97;
            32'hB0000588: data = 32'd98;
            32'hB000058C: data = 32'd99;
            32'hB0000590: data = 32'd100;
            32'hB0000594: data = 32'd101;
            32'hB0000598: data = 32'd102;
            32'hB000059C: data = 32'd103;
            32'hB00005A0: data = 32'd104;
            32'hB00005A4: data = 32'd105;
            32'hB00005A8: data = 32'd106;
            32'hB00005AC: data = 32'd107;
            32'hB00005B0: data = 32'd108;
            32'hB00005B4: data = 32'd109;
            32'hB00005B8: data = 32'd110;
            32'hB00005BC: data = 32'd111;
            32'hB00005C0: data = 32'd112;
            32'hB00005C4: data = 32'd113;
            32'hB00005C8: data = 32'd114;
            32'hB00005CC: data = 32'd115;
            32'hB00005D0: data = 32'd116;
            32'hB00005D4: data = 32'd117;
            32'hB00005D8: data = 32'd118;
            32'hB00005DC: data = 32'd119;
            32'hB00005E0: data = 32'd120;
            32'hB00005E4: data = 32'd121;
            32'hB00005E8: data = 32'd122;
            32'hB00005EC: data = 32'd123;
            32'hB00005F0: data = 32'd124;
            32'hB00005F4: data = 32'd125;
            32'hB00005F8: data = 32'd126;
            32'hB00005FC: data = 32'd127;
            32'hB0000600: data = 32'd128;
            32'hB0000604: data = 32'd129;
            32'hB0000608: data = 32'd130;
            32'hB000060C: data = 32'd131;
            32'hB0000610: data = 32'd132;
            32'hB0000614: data = 32'd133;
            32'hB0000618: data = 32'd134;
            32'hB000061C: data = 32'd135;
            32'hB0000620: data = 32'd136;
            32'hB0000624: data = 32'd137;
            32'hB0000628: data = 32'd138;
            32'hB000062C: data = 32'd139;
            32'hB0000630: data = 32'd140;
            32'hB0000634: data = 32'd141;
            32'hB0000638: data = 32'd142;
            32'hB000063C: data = 32'd143;
            32'hB0000640: data = 32'd144;
            32'hB0000644: data = 32'd145;
            32'hB0000648: data = 32'd146;
            32'hB000064C: data = 32'd147;
            32'hB0000650: data = 32'd148;
            32'hB0000654: data = 32'd149;
            32'hB0000658: data = 32'd150;
            32'hB000065C: data = 32'd151;
            32'hB0000660: data = 32'd152;
            32'hB0000664: data = 32'd153;
            32'hB0000668: data = 32'd154;
            32'hB000066C: data = 32'd155;
            32'hB0000670: data = 32'd156;
            32'hB0000674: data = 32'd157;
            32'hB0000678: data = 32'd158;
            32'hB000067C: data = 32'd159;
            32'hB0000680: data = 32'd160;
            32'hB0000684: data = 32'd161;
            32'hB0000688: data = 32'd162;
            32'hB000068C: data = 32'd163;
            32'hB0000690: data = 32'd164;
            32'hB0000694: data = 32'd165;
            32'hB0000698: data = 32'd166;
            32'hB000069C: data = 32'd167;
            32'hB00006A0: data = 32'd168;
            32'hB00006A4: data = 32'd169;
            32'hB00006A8: data = 32'd170;
            32'hB00006AC: data = 32'd171;
            32'hB00006B0: data = 32'd172;
            32'hB00006B4: data = 32'd173;
            32'hB00006B8: data = 32'd174;
            32'hB00006BC: data = 32'd175;
            32'hB00006C0: data = 32'd176;
            32'hB00006C4: data = 32'd177;
            32'hB00006C8: data = 32'd178;
            32'hB00006CC: data = 32'd179;
            32'hB00006D0: data = 32'd180;
            32'hB00006D4: data = 32'd181;
            32'hB00006D8: data = 32'd182;
            32'hB00006DC: data = 32'd183;
            32'hB00006E0: data = 32'd184;
            32'hB00006E4: data = 32'd185;
            32'hB00006E8: data = 32'd186;
            32'hB00006EC: data = 32'd187;
            32'hB00006F0: data = 32'd188;
            32'hB00006F4: data = 32'd189;
            32'hB00006F8: data = 32'd190;
            32'hB00006FC: data = 32'd191;
            32'hB0000700: data = 32'd192;
            32'hB0000704: data = 32'd193;
            32'hB0000708: data = 32'd194;
            32'hB000070C: data = 32'd195;
            32'hB0000710: data = 32'd196;
            32'hB0000714: data = 32'd197;
            32'hB0000718: data = 32'd198;
            32'hB000071C: data = 32'd199;
            32'hB0000720: data = 32'd200;
            32'hB0000724: data = 32'd201;
            32'hB0000728: data = 32'd202;
            32'hB000072C: data = 32'd203;
            32'hB0000730: data = 32'd204;
            32'hB0000734: data = 32'd205;
            32'hB0000738: data = 32'd206;
            32'hB000073C: data = 32'd207;
            32'hB0000740: data = 32'd208;
            32'hB0000744: data = 32'd209;
            32'hB0000748: data = 32'd210;
            32'hB000074C: data = 32'd211;
            32'hB0000750: data = 32'd212;
            32'hB0000754: data = 32'd213;
            32'hB0000758: data = 32'd214;
            32'hB000075C: data = 32'd215;
            32'hB0000760: data = 32'd216;
            32'hB0000764: data = 32'd217;
            32'hB0000768: data = 32'd218;
            32'hB000076C: data = 32'd219;
            32'hB0000770: data = 32'd220;
            32'hB0000774: data = 32'd221;
            32'hB0000778: data = 32'd222;
            32'hB000077C: data = 32'd223;
            32'hB0000780: data = 32'd224;
            32'hB0000784: data = 32'd225;
            32'hB0000788: data = 32'd226;
            32'hB000078C: data = 32'd227;
            32'hB0000790: data = 32'd228;
            32'hB0000794: data = 32'd229;
            32'hB0000798: data = 32'd230;
            32'hB000079C: data = 32'd231;
            32'hB00007A0: data = 32'd232;
            32'hB00007A4: data = 32'd233;
            32'hB00007A8: data = 32'd234;
            32'hB00007AC: data = 32'd235;
            32'hB00007B0: data = 32'd236;
            32'hB00007B4: data = 32'd237;
            32'hB00007B8: data = 32'd238;
            32'hB00007BC: data = 32'd239;
            32'hB00007C0: data = 32'd240;
            32'hB00007C4: data = 32'd241;
            32'hB00007C8: data = 32'd242;
            32'hB00007CC: data = 32'd243;
            32'hB00007D0: data = 32'd244;
            32'hB00007D4: data = 32'd245;
            32'hB00007D8: data = 32'd246;
            32'hB00007DC: data = 32'd247;
            32'hB00007E0: data = 32'd248;
            32'hB00007E4: data = 32'd249;
            32'hB00007E8: data = 32'd250;
            32'hB00007EC: data = 32'd251;
            32'hB00007F0: data = 32'd252;
            32'hB00007F4: data = 32'd253;
            32'hB00007F8: data = 32'd254;
            32'hB00007FC: data = 32'd255;
            32'hB0000800: data = 32'd0;
            32'hB0000804: data = 32'd1;
            32'hB0000808: data = 32'd2;
            32'hB000080C: data = 32'd3;
            32'hB0000810: data = 32'd4;
            32'hB0000814: data = 32'd5;
            32'hB0000818: data = 32'd6;
            32'hB000081C: data = 32'd7;
            32'hB0000820: data = 32'd8;
            32'hB0000824: data = 32'd9;
            32'hB0000828: data = 32'd10;
            32'hB000082C: data = 32'd11;
            32'hB0000830: data = 32'd12;
            32'hB0000834: data = 32'd13;
            32'hB0000838: data = 32'd14;
            32'hB000083C: data = 32'd15;
            32'hB0000840: data = 32'd16;
            32'hB0000844: data = 32'd17;
            32'hB0000848: data = 32'd18;
            32'hB000084C: data = 32'd19;
            32'hB0000850: data = 32'd20;
            32'hB0000854: data = 32'd21;
            32'hB0000858: data = 32'd22;
            32'hB000085C: data = 32'd23;
            32'hB0000860: data = 32'd24;
            32'hB0000864: data = 32'd25;
            32'hB0000868: data = 32'd26;
            32'hB000086C: data = 32'd27;
            32'hB0000870: data = 32'd28;
            32'hB0000874: data = 32'd29;
            32'hB0000878: data = 32'd30;
            32'hB000087C: data = 32'd31;
            32'hB0000880: data = 32'd32;
            32'hB0000884: data = 32'd33;
            32'hB0000888: data = 32'd34;
            32'hB000088C: data = 32'd35;
            32'hB0000890: data = 32'd36;
            32'hB0000894: data = 32'd37;
            32'hB0000898: data = 32'd38;
            32'hB000089C: data = 32'd39;
            32'hB00008A0: data = 32'd40;
            32'hB00008A4: data = 32'd41;
            32'hB00008A8: data = 32'd42;
            32'hB00008AC: data = 32'd43;
            32'hB00008B0: data = 32'd44;
            32'hB00008B4: data = 32'd45;
            32'hB00008B8: data = 32'd46;
            32'hB00008BC: data = 32'd47;
            32'hB00008C0: data = 32'd48;
            32'hB00008C4: data = 32'd49;
            32'hB00008C8: data = 32'd50;
            32'hB00008CC: data = 32'd51;
            32'hB00008D0: data = 32'd52;
            32'hB00008D4: data = 32'd53;
            32'hB00008D8: data = 32'd54;
            32'hB00008DC: data = 32'd55;
            32'hB00008E0: data = 32'd56;
            32'hB00008E4: data = 32'd57;
            32'hB00008E8: data = 32'd58;
            32'hB00008EC: data = 32'd59;
            32'hB00008F0: data = 32'd60;
            32'hB00008F4: data = 32'd61;
            32'hB00008F8: data = 32'd62;
            32'hB00008FC: data = 32'd63;
            32'hB0000900: data = 32'd64;
            32'hB0000904: data = 32'd65;
            32'hB0000908: data = 32'd66;
            32'hB000090C: data = 32'd67;
            32'hB0000910: data = 32'd68;
            32'hB0000914: data = 32'd69;
            32'hB0000918: data = 32'd70;
            32'hB000091C: data = 32'd71;
            32'hB0000920: data = 32'd72;
            32'hB0000924: data = 32'd73;
            32'hB0000928: data = 32'd74;
            32'hB000092C: data = 32'd75;
            32'hB0000930: data = 32'd76;
            32'hB0000934: data = 32'd77;
            32'hB0000938: data = 32'd78;
            32'hB000093C: data = 32'd79;
            32'hB0000940: data = 32'd80;
            32'hB0000944: data = 32'd81;
            32'hB0000948: data = 32'd82;
            32'hB000094C: data = 32'd83;
            32'hB0000950: data = 32'd84;
            32'hB0000954: data = 32'd85;
            32'hB0000958: data = 32'd86;
            32'hB000095C: data = 32'd87;
            32'hB0000960: data = 32'd88;
            32'hB0000964: data = 32'd89;
            32'hB0000968: data = 32'd90;
            32'hB000096C: data = 32'd91;
            32'hB0000970: data = 32'd92;
            32'hB0000974: data = 32'd93;
            32'hB0000978: data = 32'd94;
            32'hB000097C: data = 32'd95;
            32'hB0000980: data = 32'd96;
            32'hB0000984: data = 32'd97;
            32'hB0000988: data = 32'd98;
            32'hB000098C: data = 32'd99;
            32'hB0000990: data = 32'd100;
            32'hB0000994: data = 32'd101;
            32'hB0000998: data = 32'd102;
            32'hB000099C: data = 32'd103;
            32'hB00009A0: data = 32'd104;
            32'hB00009A4: data = 32'd105;
            32'hB00009A8: data = 32'd106;
            32'hB00009AC: data = 32'd107;
            32'hB00009B0: data = 32'd108;
            32'hB00009B4: data = 32'd109;
            32'hB00009B8: data = 32'd110;
            32'hB00009BC: data = 32'd111;
            32'hB00009C0: data = 32'd112;
            32'hB00009C4: data = 32'd113;
            32'hB00009C8: data = 32'd114;
            32'hB00009CC: data = 32'd115;
            32'hB00009D0: data = 32'd116;
            32'hB00009D4: data = 32'd117;
            32'hB00009D8: data = 32'd118;
            32'hB00009DC: data = 32'd119;
            32'hB00009E0: data = 32'd120;
            32'hB00009E4: data = 32'd121;
            32'hB00009E8: data = 32'd122;
            32'hB00009EC: data = 32'd123;
            32'hB00009F0: data = 32'd124;
            32'hB00009F4: data = 32'd125;
            32'hB00009F8: data = 32'd126;
            32'hB00009FC: data = 32'd127;
            32'hB0000A00: data = 32'd128;
            32'hB0000A04: data = 32'd129;
            32'hB0000A08: data = 32'd130;
            32'hB0000A0C: data = 32'd131;
            32'hB0000A10: data = 32'd132;
            32'hB0000A14: data = 32'd133;
            32'hB0000A18: data = 32'd134;
            32'hB0000A1C: data = 32'd135;
            32'hB0000A20: data = 32'd136;
            32'hB0000A24: data = 32'd137;
            32'hB0000A28: data = 32'd138;
            32'hB0000A2C: data = 32'd139;
            32'hB0000A30: data = 32'd140;
            32'hB0000A34: data = 32'd141;
            32'hB0000A38: data = 32'd142;
            32'hB0000A3C: data = 32'd143;
            32'hB0000A40: data = 32'd144;
            32'hB0000A44: data = 32'd145;
            32'hB0000A48: data = 32'd146;
            32'hB0000A4C: data = 32'd147;
            32'hB0000A50: data = 32'd148;
            32'hB0000A54: data = 32'd149;
            32'hB0000A58: data = 32'd150;
            32'hB0000A5C: data = 32'd151;
            32'hB0000A60: data = 32'd152;
            32'hB0000A64: data = 32'd153;
            32'hB0000A68: data = 32'd154;
            32'hB0000A6C: data = 32'd155;
            32'hB0000A70: data = 32'd156;
            32'hB0000A74: data = 32'd157;
            32'hB0000A78: data = 32'd158;
            32'hB0000A7C: data = 32'd159;
            32'hB0000A80: data = 32'd160;
            32'hB0000A84: data = 32'd161;
            32'hB0000A88: data = 32'd162;
            32'hB0000A8C: data = 32'd163;
            32'hB0000A90: data = 32'd164;
            32'hB0000A94: data = 32'd165;
            32'hB0000A98: data = 32'd166;
            32'hB0000A9C: data = 32'd167;
            32'hB0000AA0: data = 32'd168;
            32'hB0000AA4: data = 32'd169;
            32'hB0000AA8: data = 32'd170;
            32'hB0000AAC: data = 32'd171;
            32'hB0000AB0: data = 32'd172;
            32'hB0000AB4: data = 32'd173;
            32'hB0000AB8: data = 32'd174;
            32'hB0000ABC: data = 32'd175;
            32'hB0000AC0: data = 32'd176;
            32'hB0000AC4: data = 32'd177;
            32'hB0000AC8: data = 32'd178;
            32'hB0000ACC: data = 32'd179;
            32'hB0000AD0: data = 32'd180;
            32'hB0000AD4: data = 32'd181;
            32'hB0000AD8: data = 32'd182;
            32'hB0000ADC: data = 32'd183;
            32'hB0000AE0: data = 32'd184;
            32'hB0000AE4: data = 32'd185;
            32'hB0000AE8: data = 32'd186;
            32'hB0000AEC: data = 32'd187;
            32'hB0000AF0: data = 32'd188;
            32'hB0000AF4: data = 32'd189;
            32'hB0000AF8: data = 32'd190;
            32'hB0000AFC: data = 32'd191;
            32'hB0000B00: data = 32'd192;
            32'hB0000B04: data = 32'd193;
            32'hB0000B08: data = 32'd194;
            32'hB0000B0C: data = 32'd195;
            32'hB0000B10: data = 32'd196;
            32'hB0000B14: data = 32'd197;
            32'hB0000B18: data = 32'd198;
            32'hB0000B1C: data = 32'd199;
            32'hB0000B20: data = 32'd200;
            32'hB0000B24: data = 32'd201;
            32'hB0000B28: data = 32'd202;
            32'hB0000B2C: data = 32'd203;
            32'hB0000B30: data = 32'd204;
            32'hB0000B34: data = 32'd205;
            32'hB0000B38: data = 32'd206;
            32'hB0000B3C: data = 32'd207;
            32'hB0000B40: data = 32'd208;
            32'hB0000B44: data = 32'd209;
            32'hB0000B48: data = 32'd210;
            32'hB0000B4C: data = 32'd211;
            32'hB0000B50: data = 32'd212;
            32'hB0000B54: data = 32'd213;
            32'hB0000B58: data = 32'd214;
            32'hB0000B5C: data = 32'd215;
            32'hB0000B60: data = 32'd216;
            32'hB0000B64: data = 32'd217;
            32'hB0000B68: data = 32'd218;
            32'hB0000B6C: data = 32'd219;
            32'hB0000B70: data = 32'd220;
            32'hB0000B74: data = 32'd221;
            32'hB0000B78: data = 32'd222;
            32'hB0000B7C: data = 32'd223;
            32'hB0000B80: data = 32'd224;
            32'hB0000B84: data = 32'd225;
            32'hB0000B88: data = 32'd226;
            32'hB0000B8C: data = 32'd227;
            32'hB0000B90: data = 32'd228;
            32'hB0000B94: data = 32'd229;
            32'hB0000B98: data = 32'd230;
            32'hB0000B9C: data = 32'd231;
            32'hB0000BA0: data = 32'd232;
            32'hB0000BA4: data = 32'd233;
            32'hB0000BA8: data = 32'd234;
            32'hB0000BAC: data = 32'd235;
            32'hB0000BB0: data = 32'd236;
            32'hB0000BB4: data = 32'd237;
            32'hB0000BB8: data = 32'd238;
            32'hB0000BBC: data = 32'd239;
            32'hB0000BC0: data = 32'd240;
            32'hB0000BC4: data = 32'd241;
            32'hB0000BC8: data = 32'd242;
            32'hB0000BCC: data = 32'd243;
            32'hB0000BD0: data = 32'd244;
            32'hB0000BD4: data = 32'd245;
            32'hB0000BD8: data = 32'd246;
            32'hB0000BDC: data = 32'd247;
            32'hB0000BE0: data = 32'd248;
            32'hB0000BE4: data = 32'd249;
            32'hB0000BE8: data = 32'd250;
            32'hB0000BEC: data = 32'd251;
            32'hB0000BF0: data = 32'd252;
            32'hB0000BF4: data = 32'd253;
            32'hB0000BF8: data = 32'd254;
            32'hB0000BFC: data = 32'd255;
            32'hB0000C00: data = 32'd0;
            32'hB0000C04: data = 32'd1;
            32'hB0000C08: data = 32'd2;
            32'hB0000C0C: data = 32'd3;
            32'hB0000C10: data = 32'd4;
            32'hB0000C14: data = 32'd5;
            32'hB0000C18: data = 32'd6;
            32'hB0000C1C: data = 32'd7;
            32'hB0000C20: data = 32'd8;
            32'hB0000C24: data = 32'd9;
            32'hB0000C28: data = 32'd10;
            32'hB0000C2C: data = 32'd11;
            32'hB0000C30: data = 32'd12;
            32'hB0000C34: data = 32'd13;
            32'hB0000C38: data = 32'd14;
            32'hB0000C3C: data = 32'd15;
            32'hB0000C40: data = 32'd16;
            32'hB0000C44: data = 32'd17;
            32'hB0000C48: data = 32'd18;
            32'hB0000C4C: data = 32'd19;
            32'hB0000C50: data = 32'd20;
            32'hB0000C54: data = 32'd21;
            32'hB0000C58: data = 32'd22;
            32'hB0000C5C: data = 32'd23;
            32'hB0000C60: data = 32'd24;
            32'hB0000C64: data = 32'd25;
            32'hB0000C68: data = 32'd26;
            32'hB0000C6C: data = 32'd27;
            32'hB0000C70: data = 32'd28;
            32'hB0000C74: data = 32'd29;
            32'hB0000C78: data = 32'd30;
            32'hB0000C7C: data = 32'd31;
            32'hB0000C80: data = 32'd32;
            32'hB0000C84: data = 32'd33;
            32'hB0000C88: data = 32'd34;
            32'hB0000C8C: data = 32'd35;
            32'hB0000C90: data = 32'd36;
            32'hB0000C94: data = 32'd37;
            32'hB0000C98: data = 32'd38;
            32'hB0000C9C: data = 32'd39;
            32'hB0000CA0: data = 32'd40;
            32'hB0000CA4: data = 32'd41;
            32'hB0000CA8: data = 32'd42;
            32'hB0000CAC: data = 32'd43;
            32'hB0000CB0: data = 32'd44;
            32'hB0000CB4: data = 32'd45;
            32'hB0000CB8: data = 32'd46;
            32'hB0000CBC: data = 32'd47;
            32'hB0000CC0: data = 32'd48;
            32'hB0000CC4: data = 32'd49;
            32'hB0000CC8: data = 32'd50;
            32'hB0000CCC: data = 32'd51;
            32'hB0000CD0: data = 32'd52;
            32'hB0000CD4: data = 32'd53;
            32'hB0000CD8: data = 32'd54;
            32'hB0000CDC: data = 32'd55;
            32'hB0000CE0: data = 32'd56;
            32'hB0000CE4: data = 32'd57;
            32'hB0000CE8: data = 32'd58;
            32'hB0000CEC: data = 32'd59;
            32'hB0000CF0: data = 32'd60;
            32'hB0000CF4: data = 32'd61;
            32'hB0000CF8: data = 32'd62;
            32'hB0000CFC: data = 32'd63;
            32'hB0000D00: data = 32'd64;
            32'hB0000D04: data = 32'd65;
            32'hB0000D08: data = 32'd66;
            32'hB0000D0C: data = 32'd67;
            32'hB0000D10: data = 32'd68;
            32'hB0000D14: data = 32'd69;
            32'hB0000D18: data = 32'd70;
            32'hB0000D1C: data = 32'd71;
            32'hB0000D20: data = 32'd72;
            32'hB0000D24: data = 32'd73;
            32'hB0000D28: data = 32'd74;
            32'hB0000D2C: data = 32'd75;
            32'hB0000D30: data = 32'd76;
            32'hB0000D34: data = 32'd77;
            32'hB0000D38: data = 32'd78;
            32'hB0000D3C: data = 32'd79;
            32'hB0000D40: data = 32'd80;
            32'hB0000D44: data = 32'd81;
            32'hB0000D48: data = 32'd82;
            32'hB0000D4C: data = 32'd83;
            32'hB0000D50: data = 32'd84;
            32'hB0000D54: data = 32'd85;
            32'hB0000D58: data = 32'd86;
            32'hB0000D5C: data = 32'd87;
            32'hB0000D60: data = 32'd88;
            32'hB0000D64: data = 32'd89;
            32'hB0000D68: data = 32'd90;
            32'hB0000D6C: data = 32'd91;
            32'hB0000D70: data = 32'd92;
            32'hB0000D74: data = 32'd93;
            32'hB0000D78: data = 32'd94;
            32'hB0000D7C: data = 32'd95;
            32'hB0000D80: data = 32'd96;
            32'hB0000D84: data = 32'd97;
            32'hB0000D88: data = 32'd98;
            32'hB0000D8C: data = 32'd99;
            32'hB0000D90: data = 32'd100;
            32'hB0000D94: data = 32'd101;
            32'hB0000D98: data = 32'd102;
            32'hB0000D9C: data = 32'd103;
            32'hB0000DA0: data = 32'd104;
            32'hB0000DA4: data = 32'd105;
            32'hB0000DA8: data = 32'd106;
            32'hB0000DAC: data = 32'd107;
            32'hB0000DB0: data = 32'd108;
            32'hB0000DB4: data = 32'd109;
            32'hB0000DB8: data = 32'd110;
            32'hB0000DBC: data = 32'd111;
            32'hB0000DC0: data = 32'd112;
            32'hB0000DC4: data = 32'd113;
            32'hB0000DC8: data = 32'd114;
            32'hB0000DCC: data = 32'd115;
            32'hB0000DD0: data = 32'd116;
            32'hB0000DD4: data = 32'd117;
            32'hB0000DD8: data = 32'd118;
            32'hB0000DDC: data = 32'd119;
            32'hB0000DE0: data = 32'd120;
            32'hB0000DE4: data = 32'd121;
            32'hB0000DE8: data = 32'd122;
            32'hB0000DEC: data = 32'd123;
            32'hB0000DF0: data = 32'd124;
            32'hB0000DF4: data = 32'd125;
            32'hB0000DF8: data = 32'd126;
            32'hB0000DFC: data = 32'd127;
            32'hB0000E00: data = 32'd128;
            32'hB0000E04: data = 32'd129;
            32'hB0000E08: data = 32'd130;
            32'hB0000E0C: data = 32'd131;
            32'hB0000E10: data = 32'd132;
            32'hB0000E14: data = 32'd133;
            32'hB0000E18: data = 32'd134;
            32'hB0000E1C: data = 32'd135;
            32'hB0000E20: data = 32'd136;
            32'hB0000E24: data = 32'd137;
            32'hB0000E28: data = 32'd138;
            32'hB0000E2C: data = 32'd139;
            32'hB0000E30: data = 32'd140;
            32'hB0000E34: data = 32'd141;
            32'hB0000E38: data = 32'd142;
            32'hB0000E3C: data = 32'd143;
            32'hB0000E40: data = 32'd144;
            32'hB0000E44: data = 32'd145;
            32'hB0000E48: data = 32'd146;
            32'hB0000E4C: data = 32'd147;
            32'hB0000E50: data = 32'd148;
            32'hB0000E54: data = 32'd149;
            32'hB0000E58: data = 32'd150;
            32'hB0000E5C: data = 32'd151;
            32'hB0000E60: data = 32'd152;
            32'hB0000E64: data = 32'd153;
            32'hB0000E68: data = 32'd154;
            32'hB0000E6C: data = 32'd155;
            32'hB0000E70: data = 32'd156;
            32'hB0000E74: data = 32'd157;
            32'hB0000E78: data = 32'd158;
            32'hB0000E7C: data = 32'd159;
            32'hB0000E80: data = 32'd160;
            32'hB0000E84: data = 32'd161;
            32'hB0000E88: data = 32'd162;
            32'hB0000E8C: data = 32'd163;
            32'hB0000E90: data = 32'd164;
            32'hB0000E94: data = 32'd165;
            32'hB0000E98: data = 32'd166;
            32'hB0000E9C: data = 32'd167;
            32'hB0000EA0: data = 32'd168;
            32'hB0000EA4: data = 32'd169;
            32'hB0000EA8: data = 32'd170;
            32'hB0000EAC: data = 32'd171;
            32'hB0000EB0: data = 32'd172;
            32'hB0000EB4: data = 32'd173;
            32'hB0000EB8: data = 32'd174;
            32'hB0000EBC: data = 32'd175;
            32'hB0000EC0: data = 32'd176;
            32'hB0000EC4: data = 32'd177;
            32'hB0000EC8: data = 32'd178;
            32'hB0000ECC: data = 32'd179;
            32'hB0000ED0: data = 32'd180;
            32'hB0000ED4: data = 32'd181;
            32'hB0000ED8: data = 32'd182;
            32'hB0000EDC: data = 32'd183;
            32'hB0000EE0: data = 32'd184;
            32'hB0000EE4: data = 32'd185;
            32'hB0000EE8: data = 32'd186;
            32'hB0000EEC: data = 32'd187;
            32'hB0000EF0: data = 32'd188;
            32'hB0000EF4: data = 32'd189;
            32'hB0000EF8: data = 32'd190;
            32'hB0000EFC: data = 32'd191;
            32'hB0000F00: data = 32'd192;
            32'hB0000F04: data = 32'd193;
            32'hB0000F08: data = 32'd194;
            32'hB0000F0C: data = 32'd195;
            32'hB0000F10: data = 32'd196;
            32'hB0000F14: data = 32'd197;
            32'hB0000F18: data = 32'd198;
            32'hB0000F1C: data = 32'd199;
            32'hB0000F20: data = 32'd200;
            32'hB0000F24: data = 32'd201;
            32'hB0000F28: data = 32'd202;
            32'hB0000F2C: data = 32'd203;
            32'hB0000F30: data = 32'd204;
            32'hB0000F34: data = 32'd205;
            32'hB0000F38: data = 32'd206;
            32'hB0000F3C: data = 32'd207;
            32'hB0000F40: data = 32'd208;
            32'hB0000F44: data = 32'd209;
            32'hB0000F48: data = 32'd210;
            32'hB0000F4C: data = 32'd211;
            32'hB0000F50: data = 32'd212;
            32'hB0000F54: data = 32'd213;
            32'hB0000F58: data = 32'd214;
            32'hB0000F5C: data = 32'd215;
            32'hB0000F60: data = 32'd216;
            32'hB0000F64: data = 32'd217;
            32'hB0000F68: data = 32'd218;
            32'hB0000F6C: data = 32'd219;
            32'hB0000F70: data = 32'd220;
            32'hB0000F74: data = 32'd221;
            32'hB0000F78: data = 32'd222;
            32'hB0000F7C: data = 32'd223;
            32'hB0000F80: data = 32'd224;
            32'hB0000F84: data = 32'd225;
            32'hB0000F88: data = 32'd226;
            32'hB0000F8C: data = 32'd227;
            32'hB0000F90: data = 32'd228;
            32'hB0000F94: data = 32'd229;
            32'hB0000F98: data = 32'd230;
            32'hB0000F9C: data = 32'd231;
            32'hB0000FA0: data = 32'd232;
            32'hB0000FA4: data = 32'd233;
            32'hB0000FA8: data = 32'd234;
            32'hB0000FAC: data = 32'd235;
            32'hB0000FB0: data = 32'd236;
            32'hB0000FB4: data = 32'd237;
            32'hB0000FB8: data = 32'd238;
            32'hB0000FBC: data = 32'd239;
            32'hB0000FC0: data = 32'd240;
            32'hB0000FC4: data = 32'd241;
            32'hB0000FC8: data = 32'd242;
            32'hB0000FCC: data = 32'd243;
            32'hB0000FD0: data = 32'd244;
            32'hB0000FD4: data = 32'd245;
            32'hB0000FD8: data = 32'd246;
            32'hB0000FDC: data = 32'd247;
            32'hB0000FE0: data = 32'd248;
            32'hB0000FE4: data = 32'd249;
            32'hB0000FE8: data = 32'd250;
            32'hB0000FEC: data = 32'd251;
            32'hB0000FF0: data = 32'd252;
            32'hB0000FF4: data = 32'd253;
            32'hB0000FF8: data = 32'd254;
            32'hB0000FFC: data = 32'd255;
            32'hB0001000: data = 32'd0;
            32'hB0001004: data = 32'd1;
            32'hB0001008: data = 32'd2;
            32'hB000100C: data = 32'd3;
            32'hB0001010: data = 32'd4;
            32'hB0001014: data = 32'd5;
            32'hB0001018: data = 32'd6;
            32'hB000101C: data = 32'd7;
            32'hB0001020: data = 32'd8;
            32'hB0001024: data = 32'd9;
            32'hB0001028: data = 32'd10;
            32'hB000102C: data = 32'd11;
            32'hB0001030: data = 32'd12;
            32'hB0001034: data = 32'd13;
            32'hB0001038: data = 32'd14;
            32'hB000103C: data = 32'd15;
            32'hB0001040: data = 32'd16;
            32'hB0001044: data = 32'd17;
            32'hB0001048: data = 32'd18;
            32'hB000104C: data = 32'd19;
            32'hB0001050: data = 32'd20;
            32'hB0001054: data = 32'd21;
            32'hB0001058: data = 32'd22;
            32'hB000105C: data = 32'd23;
            32'hB0001060: data = 32'd24;
            32'hB0001064: data = 32'd25;
            32'hB0001068: data = 32'd26;
            32'hB000106C: data = 32'd27;
            32'hB0001070: data = 32'd28;
            32'hB0001074: data = 32'd29;
            32'hB0001078: data = 32'd30;
            32'hB000107C: data = 32'd31;
            32'hB0001080: data = 32'd32;
            32'hB0001084: data = 32'd33;
            32'hB0001088: data = 32'd34;
            32'hB000108C: data = 32'd35;
            32'hB0001090: data = 32'd36;
            32'hB0001094: data = 32'd37;
            32'hB0001098: data = 32'd38;
            32'hB000109C: data = 32'd39;
            32'hB00010A0: data = 32'd40;
            32'hB00010A4: data = 32'd41;
            32'hB00010A8: data = 32'd42;
            32'hB00010AC: data = 32'd43;
            32'hB00010B0: data = 32'd44;
            32'hB00010B4: data = 32'd45;
            32'hB00010B8: data = 32'd46;
            32'hB00010BC: data = 32'd47;
            32'hB00010C0: data = 32'd48;
            32'hB00010C4: data = 32'd49;
            32'hB00010C8: data = 32'd50;
            32'hB00010CC: data = 32'd51;
            32'hB00010D0: data = 32'd52;
            32'hB00010D4: data = 32'd53;
            32'hB00010D8: data = 32'd54;
            32'hB00010DC: data = 32'd55;
            32'hB00010E0: data = 32'd56;
            32'hB00010E4: data = 32'd57;
            32'hB00010E8: data = 32'd58;
            32'hB00010EC: data = 32'd59;
            32'hB00010F0: data = 32'd60;
            32'hB00010F4: data = 32'd61;
            32'hB00010F8: data = 32'd62;
            32'hB00010FC: data = 32'd63;
            32'hB0001100: data = 32'd64;
            32'hB0001104: data = 32'd65;
            32'hB0001108: data = 32'd66;
            32'hB000110C: data = 32'd67;
            32'hB0001110: data = 32'd68;
            32'hB0001114: data = 32'd69;
            32'hB0001118: data = 32'd70;
            32'hB000111C: data = 32'd71;
            32'hB0001120: data = 32'd72;
            32'hB0001124: data = 32'd73;
            32'hB0001128: data = 32'd74;
            32'hB000112C: data = 32'd75;
            32'hB0001130: data = 32'd76;
            32'hB0001134: data = 32'd77;
            32'hB0001138: data = 32'd78;
            32'hB000113C: data = 32'd79;
            32'hB0001140: data = 32'd80;
            32'hB0001144: data = 32'd81;
            32'hB0001148: data = 32'd82;
            32'hB000114C: data = 32'd83;
            32'hB0001150: data = 32'd84;
            32'hB0001154: data = 32'd85;
            32'hB0001158: data = 32'd86;
            32'hB000115C: data = 32'd87;
            32'hB0001160: data = 32'd88;
            32'hB0001164: data = 32'd89;
            32'hB0001168: data = 32'd90;
            32'hB000116C: data = 32'd91;
            32'hB0001170: data = 32'd92;
            32'hB0001174: data = 32'd93;
            32'hB0001178: data = 32'd94;
            32'hB000117C: data = 32'd95;
            32'hB0001180: data = 32'd96;
            32'hB0001184: data = 32'd97;
            32'hB0001188: data = 32'd98;
            32'hB000118C: data = 32'd99;
            32'hB0001190: data = 32'd100;
            32'hB0001194: data = 32'd101;
            32'hB0001198: data = 32'd102;
            32'hB000119C: data = 32'd103;
            32'hB00011A0: data = 32'd104;
            32'hB00011A4: data = 32'd105;
            32'hB00011A8: data = 32'd106;
            32'hB00011AC: data = 32'd107;
            32'hB00011B0: data = 32'd108;
            32'hB00011B4: data = 32'd109;
            32'hB00011B8: data = 32'd110;
            32'hB00011BC: data = 32'd111;
            32'hB00011C0: data = 32'd112;
            32'hB00011C4: data = 32'd113;
            32'hB00011C8: data = 32'd114;
            32'hB00011CC: data = 32'd115;
            32'hB00011D0: data = 32'd116;
            32'hB00011D4: data = 32'd117;
            32'hB00011D8: data = 32'd118;
            32'hB00011DC: data = 32'd119;
            32'hB00011E0: data = 32'd120;
            32'hB00011E4: data = 32'd121;
            32'hB00011E8: data = 32'd122;
            32'hB00011EC: data = 32'd123;
            32'hB00011F0: data = 32'd124;
            32'hB00011F4: data = 32'd125;
            32'hB00011F8: data = 32'd126;
            32'hB00011FC: data = 32'd127;
            32'hB0001200: data = 32'd128;
            32'hB0001204: data = 32'd129;
            32'hB0001208: data = 32'd130;
            32'hB000120C: data = 32'd131;
            32'hB0001210: data = 32'd132;
            32'hB0001214: data = 32'd133;
            32'hB0001218: data = 32'd134;
            32'hB000121C: data = 32'd135;
            32'hB0001220: data = 32'd136;
            32'hB0001224: data = 32'd137;
            32'hB0001228: data = 32'd138;
            32'hB000122C: data = 32'd139;
            32'hB0001230: data = 32'd140;
            32'hB0001234: data = 32'd141;
            32'hB0001238: data = 32'd142;
            32'hB000123C: data = 32'd143;
            32'hB0001240: data = 32'd144;
            32'hB0001244: data = 32'd145;
            32'hB0001248: data = 32'd146;
            32'hB000124C: data = 32'd147;
            32'hB0001250: data = 32'd148;
            32'hB0001254: data = 32'd149;
            32'hB0001258: data = 32'd150;
            32'hB000125C: data = 32'd151;
            32'hB0001260: data = 32'd152;
            32'hB0001264: data = 32'd153;
            32'hB0001268: data = 32'd154;
            32'hB000126C: data = 32'd155;
            32'hB0001270: data = 32'd156;
            32'hB0001274: data = 32'd157;
            32'hB0001278: data = 32'd158;
            32'hB000127C: data = 32'd159;
            32'hB0001280: data = 32'd160;
            32'hB0001284: data = 32'd161;
            32'hB0001288: data = 32'd162;
            32'hB000128C: data = 32'd163;
            32'hB0001290: data = 32'd164;
            32'hB0001294: data = 32'd165;
            32'hB0001298: data = 32'd166;
            32'hB000129C: data = 32'd167;
            32'hB00012A0: data = 32'd168;
            32'hB00012A4: data = 32'd169;
            32'hB00012A8: data = 32'd170;
            32'hB00012AC: data = 32'd171;
            32'hB00012B0: data = 32'd172;
            32'hB00012B4: data = 32'd173;
            32'hB00012B8: data = 32'd174;
            32'hB00012BC: data = 32'd175;
            32'hB00012C0: data = 32'd176;
            32'hB00012C4: data = 32'd177;
            32'hB00012C8: data = 32'd178;
            32'hB00012CC: data = 32'd179;
            32'hB00012D0: data = 32'd180;
            32'hB00012D4: data = 32'd181;
            32'hB00012D8: data = 32'd182;
            32'hB00012DC: data = 32'd183;
            32'hB00012E0: data = 32'd184;
            32'hB00012E4: data = 32'd185;
            32'hB00012E8: data = 32'd186;
            32'hB00012EC: data = 32'd187;
            32'hB00012F0: data = 32'd188;
            32'hB00012F4: data = 32'd189;
            32'hB00012F8: data = 32'd190;
            32'hB00012FC: data = 32'd191;
            32'hB0001300: data = 32'd192;
            32'hB0001304: data = 32'd193;
            32'hB0001308: data = 32'd194;
            32'hB000130C: data = 32'd195;
            32'hB0001310: data = 32'd196;
            32'hB0001314: data = 32'd197;
            32'hB0001318: data = 32'd198;
            32'hB000131C: data = 32'd199;
            32'hB0001320: data = 32'd200;
            32'hB0001324: data = 32'd201;
            32'hB0001328: data = 32'd202;
            32'hB000132C: data = 32'd203;
            32'hB0001330: data = 32'd204;
            32'hB0001334: data = 32'd205;
            32'hB0001338: data = 32'd206;
            32'hB000133C: data = 32'd207;
            32'hB0001340: data = 32'd208;
            32'hB0001344: data = 32'd209;
            32'hB0001348: data = 32'd210;
            32'hB000134C: data = 32'd211;
            32'hB0001350: data = 32'd212;
            32'hB0001354: data = 32'd213;
            32'hB0001358: data = 32'd214;
            32'hB000135C: data = 32'd215;
            32'hB0001360: data = 32'd216;
            32'hB0001364: data = 32'd217;
            32'hB0001368: data = 32'd218;
            32'hB000136C: data = 32'd219;
            32'hB0001370: data = 32'd220;
            32'hB0001374: data = 32'd221;
            32'hB0001378: data = 32'd222;
            32'hB000137C: data = 32'd223;
            32'hB0001380: data = 32'd224;
            32'hB0001384: data = 32'd225;
            32'hB0001388: data = 32'd226;
            32'hB000138C: data = 32'd227;
            32'hB0001390: data = 32'd228;
            32'hB0001394: data = 32'd229;
            32'hB0001398: data = 32'd230;
            32'hB000139C: data = 32'd231;
            32'hB00013A0: data = 32'd232;
            32'hB00013A4: data = 32'd233;
            32'hB00013A8: data = 32'd234;
            32'hB00013AC: data = 32'd235;
            32'hB00013B0: data = 32'd236;
            32'hB00013B4: data = 32'd237;
            32'hB00013B8: data = 32'd238;
            32'hB00013BC: data = 32'd239;
            32'hB00013C0: data = 32'd240;
            32'hB00013C4: data = 32'd241;
            32'hB00013C8: data = 32'd242;
            32'hB00013CC: data = 32'd243;
            32'hB00013D0: data = 32'd244;
            32'hB00013D4: data = 32'd245;
            32'hB00013D8: data = 32'd246;
            32'hB00013DC: data = 32'd247;
            32'hB00013E0: data = 32'd248;
            32'hB00013E4: data = 32'd249;
            32'hB00013E8: data = 32'd250;
            32'hB00013EC: data = 32'd251;
            32'hB00013F0: data = 32'd252;
            32'hB00013F4: data = 32'd253;
            32'hB00013F8: data = 32'd254;
            32'hB00013FC: data = 32'd255;
            32'hB0001400: data = 32'd0;
            32'hB0001404: data = 32'd1;
            32'hB0001408: data = 32'd2;
            32'hB000140C: data = 32'd3;
            32'hB0001410: data = 32'd4;
            32'hB0001414: data = 32'd5;
            32'hB0001418: data = 32'd6;
            32'hB000141C: data = 32'd7;
            32'hB0001420: data = 32'd8;
            32'hB0001424: data = 32'd9;
            32'hB0001428: data = 32'd10;
            32'hB000142C: data = 32'd11;
            32'hB0001430: data = 32'd12;
            32'hB0001434: data = 32'd13;
            32'hB0001438: data = 32'd14;
            32'hB000143C: data = 32'd15;
            32'hB0001440: data = 32'd16;
            32'hB0001444: data = 32'd17;
            32'hB0001448: data = 32'd18;
            32'hB000144C: data = 32'd19;
            32'hB0001450: data = 32'd20;
            32'hB0001454: data = 32'd21;
            32'hB0001458: data = 32'd22;
            32'hB000145C: data = 32'd23;
            32'hB0001460: data = 32'd24;
            32'hB0001464: data = 32'd25;
            32'hB0001468: data = 32'd26;
            32'hB000146C: data = 32'd27;
            32'hB0001470: data = 32'd28;
            32'hB0001474: data = 32'd29;
            32'hB0001478: data = 32'd30;
            32'hB000147C: data = 32'd31;
            32'hB0001480: data = 32'd32;
            32'hB0001484: data = 32'd33;
            32'hB0001488: data = 32'd34;
            32'hB000148C: data = 32'd35;
            32'hB0001490: data = 32'd36;
            32'hB0001494: data = 32'd37;
            32'hB0001498: data = 32'd38;
            32'hB000149C: data = 32'd39;
            32'hB00014A0: data = 32'd40;
            32'hB00014A4: data = 32'd41;
            32'hB00014A8: data = 32'd42;
            32'hB00014AC: data = 32'd43;
            32'hB00014B0: data = 32'd44;
            32'hB00014B4: data = 32'd45;
            32'hB00014B8: data = 32'd46;
            32'hB00014BC: data = 32'd47;
            32'hB00014C0: data = 32'd48;
            32'hB00014C4: data = 32'd49;
            32'hB00014C8: data = 32'd50;
            32'hB00014CC: data = 32'd51;
            32'hB00014D0: data = 32'd52;
            32'hB00014D4: data = 32'd53;
            32'hB00014D8: data = 32'd54;
            32'hB00014DC: data = 32'd55;
            32'hB00014E0: data = 32'd56;
            32'hB00014E4: data = 32'd57;
            32'hB00014E8: data = 32'd58;
            32'hB00014EC: data = 32'd59;
            32'hB00014F0: data = 32'd60;
            32'hB00014F4: data = 32'd61;
            32'hB00014F8: data = 32'd62;
            32'hB00014FC: data = 32'd63;
            32'hB0001500: data = 32'd64;
            32'hB0001504: data = 32'd65;
            32'hB0001508: data = 32'd66;
            32'hB000150C: data = 32'd67;
            32'hB0001510: data = 32'd68;
            32'hB0001514: data = 32'd69;
            32'hB0001518: data = 32'd70;
            32'hB000151C: data = 32'd71;
            32'hB0001520: data = 32'd72;
            32'hB0001524: data = 32'd73;
            32'hB0001528: data = 32'd74;
            32'hB000152C: data = 32'd75;
            32'hB0001530: data = 32'd76;
            32'hB0001534: data = 32'd77;
            32'hB0001538: data = 32'd78;
            32'hB000153C: data = 32'd79;
            32'hB0001540: data = 32'd80;
            32'hB0001544: data = 32'd81;
            32'hB0001548: data = 32'd82;
            32'hB000154C: data = 32'd83;
            32'hB0001550: data = 32'd84;
            32'hB0001554: data = 32'd85;
            32'hB0001558: data = 32'd86;
            32'hB000155C: data = 32'd87;
            32'hB0001560: data = 32'd88;
            32'hB0001564: data = 32'd89;
            32'hB0001568: data = 32'd90;
            32'hB000156C: data = 32'd91;
            32'hB0001570: data = 32'd92;
            32'hB0001574: data = 32'd93;
            32'hB0001578: data = 32'd94;
            32'hB000157C: data = 32'd95;
            32'hB0001580: data = 32'd96;
            32'hB0001584: data = 32'd97;
            32'hB0001588: data = 32'd98;
            32'hB000158C: data = 32'd99;
            32'hB0001590: data = 32'd100;
            32'hB0001594: data = 32'd101;
            32'hB0001598: data = 32'd102;
            32'hB000159C: data = 32'd103;
            32'hB00015A0: data = 32'd104;
            32'hB00015A4: data = 32'd105;
            32'hB00015A8: data = 32'd106;
            32'hB00015AC: data = 32'd107;
            32'hB00015B0: data = 32'd108;
            32'hB00015B4: data = 32'd109;
            32'hB00015B8: data = 32'd110;
            32'hB00015BC: data = 32'd111;
            32'hB00015C0: data = 32'd112;
            32'hB00015C4: data = 32'd113;
            32'hB00015C8: data = 32'd114;
            32'hB00015CC: data = 32'd115;
            32'hB00015D0: data = 32'd116;
            32'hB00015D4: data = 32'd117;
            32'hB00015D8: data = 32'd118;
            32'hB00015DC: data = 32'd119;
            32'hB00015E0: data = 32'd120;
            32'hB00015E4: data = 32'd121;
            32'hB00015E8: data = 32'd122;
            32'hB00015EC: data = 32'd123;
            32'hB00015F0: data = 32'd124;
            32'hB00015F4: data = 32'd125;
            32'hB00015F8: data = 32'd126;
            32'hB00015FC: data = 32'd127;
            32'hB0001600: data = 32'd128;
            32'hB0001604: data = 32'd129;
            32'hB0001608: data = 32'd130;
            32'hB000160C: data = 32'd131;
            32'hB0001610: data = 32'd132;
            32'hB0001614: data = 32'd133;
            32'hB0001618: data = 32'd134;
            32'hB000161C: data = 32'd135;
            32'hB0001620: data = 32'd136;
            32'hB0001624: data = 32'd137;
            32'hB0001628: data = 32'd138;
            32'hB000162C: data = 32'd139;
            32'hB0001630: data = 32'd140;
            32'hB0001634: data = 32'd141;
            32'hB0001638: data = 32'd142;
            32'hB000163C: data = 32'd143;
            32'hB0001640: data = 32'd144;
            32'hB0001644: data = 32'd145;
            32'hB0001648: data = 32'd146;
            32'hB000164C: data = 32'd147;
            32'hB0001650: data = 32'd148;
            32'hB0001654: data = 32'd149;
            32'hB0001658: data = 32'd150;
            32'hB000165C: data = 32'd151;
            32'hB0001660: data = 32'd152;
            32'hB0001664: data = 32'd153;
            32'hB0001668: data = 32'd154;
            32'hB000166C: data = 32'd155;
            32'hB0001670: data = 32'd156;
            32'hB0001674: data = 32'd157;
            32'hB0001678: data = 32'd158;
            32'hB000167C: data = 32'd159;
            32'hB0001680: data = 32'd160;
            32'hB0001684: data = 32'd161;
            32'hB0001688: data = 32'd162;
            32'hB000168C: data = 32'd163;
            32'hB0001690: data = 32'd164;
            32'hB0001694: data = 32'd165;
            32'hB0001698: data = 32'd166;
            32'hB000169C: data = 32'd167;
            32'hB00016A0: data = 32'd168;
            32'hB00016A4: data = 32'd169;
            32'hB00016A8: data = 32'd170;
            32'hB00016AC: data = 32'd171;
            32'hB00016B0: data = 32'd172;
            32'hB00016B4: data = 32'd173;
            32'hB00016B8: data = 32'd174;
            32'hB00016BC: data = 32'd175;
            32'hB00016C0: data = 32'd176;
            32'hB00016C4: data = 32'd177;
            32'hB00016C8: data = 32'd178;
            32'hB00016CC: data = 32'd179;
            32'hB00016D0: data = 32'd180;
            32'hB00016D4: data = 32'd181;
            32'hB00016D8: data = 32'd182;
            32'hB00016DC: data = 32'd183;
            32'hB00016E0: data = 32'd184;
            32'hB00016E4: data = 32'd185;
            32'hB00016E8: data = 32'd186;
            32'hB00016EC: data = 32'd187;
            32'hB00016F0: data = 32'd188;
            32'hB00016F4: data = 32'd189;
            32'hB00016F8: data = 32'd190;
            32'hB00016FC: data = 32'd191;
            32'hB0001700: data = 32'd192;
            32'hB0001704: data = 32'd193;
            32'hB0001708: data = 32'd194;
            32'hB000170C: data = 32'd195;
            32'hB0001710: data = 32'd196;
            32'hB0001714: data = 32'd197;
            32'hB0001718: data = 32'd198;
            32'hB000171C: data = 32'd199;
            32'hB0001720: data = 32'd200;
            32'hB0001724: data = 32'd201;
            32'hB0001728: data = 32'd202;
            32'hB000172C: data = 32'd203;
            32'hB0001730: data = 32'd204;
            32'hB0001734: data = 32'd205;
            32'hB0001738: data = 32'd206;
            32'hB000173C: data = 32'd207;
            32'hB0001740: data = 32'd208;
            32'hB0001744: data = 32'd209;
            32'hB0001748: data = 32'd210;
            32'hB000174C: data = 32'd211;
            32'hB0001750: data = 32'd212;
            32'hB0001754: data = 32'd213;
            32'hB0001758: data = 32'd214;
            32'hB000175C: data = 32'd215;
            32'hB0001760: data = 32'd216;
            32'hB0001764: data = 32'd217;
            32'hB0001768: data = 32'd218;
            32'hB000176C: data = 32'd219;
            32'hB0001770: data = 32'd220;
            32'hB0001774: data = 32'd221;
            32'hB0001778: data = 32'd222;
            32'hB000177C: data = 32'd223;
            32'hB0001780: data = 32'd224;
            32'hB0001784: data = 32'd225;
            32'hB0001788: data = 32'd226;
            32'hB000178C: data = 32'd227;
            32'hB0001790: data = 32'd228;
            32'hB0001794: data = 32'd229;
            32'hB0001798: data = 32'd230;
            32'hB000179C: data = 32'd231;
            32'hB00017A0: data = 32'd232;
            32'hB00017A4: data = 32'd233;
            32'hB00017A8: data = 32'd234;
            32'hB00017AC: data = 32'd235;
            32'hB00017B0: data = 32'd236;
            32'hB00017B4: data = 32'd237;
            32'hB00017B8: data = 32'd238;
            32'hB00017BC: data = 32'd239;
            32'hB00017C0: data = 32'd240;
            32'hB00017C4: data = 32'd241;
            32'hB00017C8: data = 32'd242;
            32'hB00017CC: data = 32'd243;
            32'hB00017D0: data = 32'd244;
            32'hB00017D4: data = 32'd245;
            32'hB00017D8: data = 32'd246;
            32'hB00017DC: data = 32'd247;
            32'hB00017E0: data = 32'd248;
            32'hB00017E4: data = 32'd249;
            32'hB00017E8: data = 32'd250;
            32'hB00017EC: data = 32'd251;
            32'hB00017F0: data = 32'd252;
            32'hB00017F4: data = 32'd253;
            32'hB00017F8: data = 32'd254;
            32'hB00017FC: data = 32'd255;
            32'hB0001800: data = 32'd0;
            32'hB0001804: data = 32'd1;
            32'hB0001808: data = 32'd2;
            32'hB000180C: data = 32'd3;
            32'hB0001810: data = 32'd4;
            32'hB0001814: data = 32'd5;
            32'hB0001818: data = 32'd6;
            32'hB000181C: data = 32'd7;
            32'hB0001820: data = 32'd8;
            32'hB0001824: data = 32'd9;
            32'hB0001828: data = 32'd10;
            32'hB000182C: data = 32'd11;
            32'hB0001830: data = 32'd12;
            32'hB0001834: data = 32'd13;
            32'hB0001838: data = 32'd14;
            32'hB000183C: data = 32'd15;
            32'hB0001840: data = 32'd16;
            32'hB0001844: data = 32'd17;
            32'hB0001848: data = 32'd18;
            32'hB000184C: data = 32'd19;
            32'hB0001850: data = 32'd20;
            32'hB0001854: data = 32'd21;
            32'hB0001858: data = 32'd22;
            32'hB000185C: data = 32'd23;
            32'hB0001860: data = 32'd24;
            32'hB0001864: data = 32'd25;
            32'hB0001868: data = 32'd26;
            32'hB000186C: data = 32'd27;
            32'hB0001870: data = 32'd28;
            32'hB0001874: data = 32'd29;
            32'hB0001878: data = 32'd30;
            32'hB000187C: data = 32'd31;
            32'hB0001880: data = 32'd32;
            32'hB0001884: data = 32'd33;
            32'hB0001888: data = 32'd34;
            32'hB000188C: data = 32'd35;
            32'hB0001890: data = 32'd36;
            32'hB0001894: data = 32'd37;
            32'hB0001898: data = 32'd38;
            32'hB000189C: data = 32'd39;
            32'hB00018A0: data = 32'd40;
            32'hB00018A4: data = 32'd41;
            32'hB00018A8: data = 32'd42;
            32'hB00018AC: data = 32'd43;
            32'hB00018B0: data = 32'd44;
            32'hB00018B4: data = 32'd45;
            32'hB00018B8: data = 32'd46;
            32'hB00018BC: data = 32'd47;
            32'hB00018C0: data = 32'd48;
            32'hB00018C4: data = 32'd49;
            32'hB00018C8: data = 32'd50;
            32'hB00018CC: data = 32'd51;
            32'hB00018D0: data = 32'd52;
            32'hB00018D4: data = 32'd53;
            32'hB00018D8: data = 32'd54;
            32'hB00018DC: data = 32'd55;
            32'hB00018E0: data = 32'd56;
            32'hB00018E4: data = 32'd57;
            32'hB00018E8: data = 32'd58;
            32'hB00018EC: data = 32'd59;
            32'hB00018F0: data = 32'd60;
            32'hB00018F4: data = 32'd61;
            32'hB00018F8: data = 32'd62;
            32'hB00018FC: data = 32'd63;
            32'hB0001900: data = 32'd64;
            32'hB0001904: data = 32'd65;
            32'hB0001908: data = 32'd66;
            32'hB000190C: data = 32'd67;
            32'hB0001910: data = 32'd68;
            32'hB0001914: data = 32'd69;
            32'hB0001918: data = 32'd70;
            32'hB000191C: data = 32'd71;
            32'hB0001920: data = 32'd72;
            32'hB0001924: data = 32'd73;
            32'hB0001928: data = 32'd74;
            32'hB000192C: data = 32'd75;
            32'hB0001930: data = 32'd76;
            32'hB0001934: data = 32'd77;
            32'hB0001938: data = 32'd78;
            32'hB000193C: data = 32'd79;
            32'hB0001940: data = 32'd80;
            32'hB0001944: data = 32'd81;
            32'hB0001948: data = 32'd82;
            32'hB000194C: data = 32'd83;
            32'hB0001950: data = 32'd84;
            32'hB0001954: data = 32'd85;
            32'hB0001958: data = 32'd86;
            32'hB000195C: data = 32'd87;
            32'hB0001960: data = 32'd88;
            32'hB0001964: data = 32'd89;
            32'hB0001968: data = 32'd90;
            32'hB000196C: data = 32'd91;
            32'hB0001970: data = 32'd92;
            32'hB0001974: data = 32'd93;
            32'hB0001978: data = 32'd94;
            32'hB000197C: data = 32'd95;
            32'hB0001980: data = 32'd96;
            32'hB0001984: data = 32'd97;
            32'hB0001988: data = 32'd98;
            32'hB000198C: data = 32'd99;
            32'hB0001990: data = 32'd100;
            32'hB0001994: data = 32'd101;
            32'hB0001998: data = 32'd102;
            32'hB000199C: data = 32'd103;
            32'hB00019A0: data = 32'd104;
            32'hB00019A4: data = 32'd105;
            32'hB00019A8: data = 32'd106;
            32'hB00019AC: data = 32'd107;
            32'hB00019B0: data = 32'd108;
            32'hB00019B4: data = 32'd109;
            32'hB00019B8: data = 32'd110;
            32'hB00019BC: data = 32'd111;
            32'hB00019C0: data = 32'd112;
            32'hB00019C4: data = 32'd113;
            32'hB00019C8: data = 32'd114;
            32'hB00019CC: data = 32'd115;
            32'hB00019D0: data = 32'd116;
            32'hB00019D4: data = 32'd117;
            32'hB00019D8: data = 32'd118;
            32'hB00019DC: data = 32'd119;
            32'hB00019E0: data = 32'd120;
            32'hB00019E4: data = 32'd121;
            32'hB00019E8: data = 32'd122;
            32'hB00019EC: data = 32'd123;
            32'hB00019F0: data = 32'd124;
            32'hB00019F4: data = 32'd125;
            32'hB00019F8: data = 32'd126;
            32'hB00019FC: data = 32'd127;
            32'hB0001A00: data = 32'd128;
            32'hB0001A04: data = 32'd129;
            32'hB0001A08: data = 32'd130;
            32'hB0001A0C: data = 32'd131;
            32'hB0001A10: data = 32'd132;
            32'hB0001A14: data = 32'd133;
            32'hB0001A18: data = 32'd134;
            32'hB0001A1C: data = 32'd135;
            32'hB0001A20: data = 32'd136;
            32'hB0001A24: data = 32'd137;
            32'hB0001A28: data = 32'd138;
            32'hB0001A2C: data = 32'd139;
            32'hB0001A30: data = 32'd140;
            32'hB0001A34: data = 32'd141;
            32'hB0001A38: data = 32'd142;
            32'hB0001A3C: data = 32'd143;
            32'hB0001A40: data = 32'd144;
            32'hB0001A44: data = 32'd145;
            32'hB0001A48: data = 32'd146;
            32'hB0001A4C: data = 32'd147;
            32'hB0001A50: data = 32'd148;
            32'hB0001A54: data = 32'd149;
            32'hB0001A58: data = 32'd150;
            32'hB0001A5C: data = 32'd151;
            32'hB0001A60: data = 32'd152;
            32'hB0001A64: data = 32'd153;
            32'hB0001A68: data = 32'd154;
            32'hB0001A6C: data = 32'd155;
            32'hB0001A70: data = 32'd156;
            32'hB0001A74: data = 32'd157;
            32'hB0001A78: data = 32'd158;
            32'hB0001A7C: data = 32'd159;
            32'hB0001A80: data = 32'd160;
            32'hB0001A84: data = 32'd161;
            32'hB0001A88: data = 32'd162;
            32'hB0001A8C: data = 32'd163;
            32'hB0001A90: data = 32'd164;
            32'hB0001A94: data = 32'd165;
            32'hB0001A98: data = 32'd166;
            32'hB0001A9C: data = 32'd167;
            32'hB0001AA0: data = 32'd168;
            32'hB0001AA4: data = 32'd169;
            32'hB0001AA8: data = 32'd170;
            32'hB0001AAC: data = 32'd171;
            32'hB0001AB0: data = 32'd172;
            32'hB0001AB4: data = 32'd173;
            32'hB0001AB8: data = 32'd174;
            32'hB0001ABC: data = 32'd175;
            32'hB0001AC0: data = 32'd176;
            32'hB0001AC4: data = 32'd177;
            32'hB0001AC8: data = 32'd178;
            32'hB0001ACC: data = 32'd179;
            32'hB0001AD0: data = 32'd180;
            32'hB0001AD4: data = 32'd181;
            32'hB0001AD8: data = 32'd182;
            32'hB0001ADC: data = 32'd183;
            32'hB0001AE0: data = 32'd184;
            32'hB0001AE4: data = 32'd185;
            32'hB0001AE8: data = 32'd186;
            32'hB0001AEC: data = 32'd187;
            32'hB0001AF0: data = 32'd188;
            32'hB0001AF4: data = 32'd189;
            32'hB0001AF8: data = 32'd190;
            32'hB0001AFC: data = 32'd191;
            32'hB0001B00: data = 32'd192;
            32'hB0001B04: data = 32'd193;
            32'hB0001B08: data = 32'd194;
            32'hB0001B0C: data = 32'd195;
            32'hB0001B10: data = 32'd196;
            32'hB0001B14: data = 32'd197;
            32'hB0001B18: data = 32'd198;
            32'hB0001B1C: data = 32'd199;
            32'hB0001B20: data = 32'd200;
            32'hB0001B24: data = 32'd201;
            32'hB0001B28: data = 32'd202;
            32'hB0001B2C: data = 32'd203;
            32'hB0001B30: data = 32'd204;
            32'hB0001B34: data = 32'd205;
            32'hB0001B38: data = 32'd206;
            32'hB0001B3C: data = 32'd207;
            32'hB0001B40: data = 32'd208;
            32'hB0001B44: data = 32'd209;
            32'hB0001B48: data = 32'd210;
            32'hB0001B4C: data = 32'd211;
            32'hB0001B50: data = 32'd212;
            32'hB0001B54: data = 32'd213;
            32'hB0001B58: data = 32'd214;
            32'hB0001B5C: data = 32'd215;
            32'hB0001B60: data = 32'd216;
            32'hB0001B64: data = 32'd217;
            32'hB0001B68: data = 32'd218;
            32'hB0001B6C: data = 32'd219;
            32'hB0001B70: data = 32'd220;
            32'hB0001B74: data = 32'd221;
            32'hB0001B78: data = 32'd222;
            32'hB0001B7C: data = 32'd223;
            32'hB0001B80: data = 32'd224;
            32'hB0001B84: data = 32'd225;
            32'hB0001B88: data = 32'd226;
            32'hB0001B8C: data = 32'd227;
            32'hB0001B90: data = 32'd228;
            32'hB0001B94: data = 32'd229;
            32'hB0001B98: data = 32'd230;
            32'hB0001B9C: data = 32'd231;
            32'hB0001BA0: data = 32'd232;
            32'hB0001BA4: data = 32'd233;
            32'hB0001BA8: data = 32'd234;
            32'hB0001BAC: data = 32'd235;
            32'hB0001BB0: data = 32'd236;
            32'hB0001BB4: data = 32'd237;
            32'hB0001BB8: data = 32'd238;
            32'hB0001BBC: data = 32'd239;
            32'hB0001BC0: data = 32'd240;
            32'hB0001BC4: data = 32'd241;
            32'hB0001BC8: data = 32'd242;
            32'hB0001BCC: data = 32'd243;
            32'hB0001BD0: data = 32'd244;
            32'hB0001BD4: data = 32'd245;
            32'hB0001BD8: data = 32'd246;
            32'hB0001BDC: data = 32'd247;
            32'hB0001BE0: data = 32'd248;
            32'hB0001BE4: data = 32'd249;
            32'hB0001BE8: data = 32'd250;
            32'hB0001BEC: data = 32'd251;
            32'hB0001BF0: data = 32'd252;
            32'hB0001BF4: data = 32'd253;
            32'hB0001BF8: data = 32'd254;
            32'hB0001BFC: data = 32'd255;
            32'hB0001C00: data = 32'd0;
            32'hB0001C04: data = 32'd1;
            32'hB0001C08: data = 32'd2;
            32'hB0001C0C: data = 32'd3;
            32'hB0001C10: data = 32'd4;
            32'hB0001C14: data = 32'd5;
            32'hB0001C18: data = 32'd6;
            32'hB0001C1C: data = 32'd7;
            32'hB0001C20: data = 32'd8;
            32'hB0001C24: data = 32'd9;
            32'hB0001C28: data = 32'd10;
            32'hB0001C2C: data = 32'd11;
            32'hB0001C30: data = 32'd12;
            32'hB0001C34: data = 32'd13;
            32'hB0001C38: data = 32'd14;
            32'hB0001C3C: data = 32'd15;
            32'hB0001C40: data = 32'd16;
            32'hB0001C44: data = 32'd17;
            32'hB0001C48: data = 32'd18;
            32'hB0001C4C: data = 32'd19;
            32'hB0001C50: data = 32'd20;
            32'hB0001C54: data = 32'd21;
            32'hB0001C58: data = 32'd22;
            32'hB0001C5C: data = 32'd23;
            32'hB0001C60: data = 32'd24;
            32'hB0001C64: data = 32'd25;
            32'hB0001C68: data = 32'd26;
            32'hB0001C6C: data = 32'd27;
            32'hB0001C70: data = 32'd28;
            32'hB0001C74: data = 32'd29;
            32'hB0001C78: data = 32'd30;
            32'hB0001C7C: data = 32'd31;
            32'hB0001C80: data = 32'd32;
            32'hB0001C84: data = 32'd33;
            32'hB0001C88: data = 32'd34;
            32'hB0001C8C: data = 32'd35;
            32'hB0001C90: data = 32'd36;
            32'hB0001C94: data = 32'd37;
            32'hB0001C98: data = 32'd38;
            32'hB0001C9C: data = 32'd39;
            32'hB0001CA0: data = 32'd40;
            32'hB0001CA4: data = 32'd41;
            32'hB0001CA8: data = 32'd42;
            32'hB0001CAC: data = 32'd43;
            32'hB0001CB0: data = 32'd44;
            32'hB0001CB4: data = 32'd45;
            32'hB0001CB8: data = 32'd46;
            32'hB0001CBC: data = 32'd47;
            32'hB0001CC0: data = 32'd48;
            32'hB0001CC4: data = 32'd49;
            32'hB0001CC8: data = 32'd50;
            32'hB0001CCC: data = 32'd51;
            32'hB0001CD0: data = 32'd52;
            32'hB0001CD4: data = 32'd53;
            32'hB0001CD8: data = 32'd54;
            32'hB0001CDC: data = 32'd55;
            32'hB0001CE0: data = 32'd56;
            32'hB0001CE4: data = 32'd57;
            32'hB0001CE8: data = 32'd58;
            32'hB0001CEC: data = 32'd59;
            32'hB0001CF0: data = 32'd60;
            32'hB0001CF4: data = 32'd61;
            32'hB0001CF8: data = 32'd62;
            32'hB0001CFC: data = 32'd63;
            32'hB0001D00: data = 32'd64;
            32'hB0001D04: data = 32'd65;
            32'hB0001D08: data = 32'd66;
            32'hB0001D0C: data = 32'd67;
            32'hB0001D10: data = 32'd68;
            32'hB0001D14: data = 32'd69;
            32'hB0001D18: data = 32'd70;
            32'hB0001D1C: data = 32'd71;
            32'hB0001D20: data = 32'd72;
            32'hB0001D24: data = 32'd73;
            32'hB0001D28: data = 32'd74;
            32'hB0001D2C: data = 32'd75;
            32'hB0001D30: data = 32'd76;
            32'hB0001D34: data = 32'd77;
            32'hB0001D38: data = 32'd78;
            32'hB0001D3C: data = 32'd79;
            32'hB0001D40: data = 32'd80;
            32'hB0001D44: data = 32'd81;
            32'hB0001D48: data = 32'd82;
            32'hB0001D4C: data = 32'd83;
            32'hB0001D50: data = 32'd84;
            32'hB0001D54: data = 32'd85;
            32'hB0001D58: data = 32'd86;
            32'hB0001D5C: data = 32'd87;
            32'hB0001D60: data = 32'd88;
            32'hB0001D64: data = 32'd89;
            32'hB0001D68: data = 32'd90;
            32'hB0001D6C: data = 32'd91;
            32'hB0001D70: data = 32'd92;
            32'hB0001D74: data = 32'd93;
            32'hB0001D78: data = 32'd94;
            32'hB0001D7C: data = 32'd95;
            32'hB0001D80: data = 32'd96;
            32'hB0001D84: data = 32'd97;
            32'hB0001D88: data = 32'd98;
            32'hB0001D8C: data = 32'd99;
            32'hB0001D90: data = 32'd100;
            32'hB0001D94: data = 32'd101;
            32'hB0001D98: data = 32'd102;
            32'hB0001D9C: data = 32'd103;
            32'hB0001DA0: data = 32'd104;
            32'hB0001DA4: data = 32'd105;
            32'hB0001DA8: data = 32'd106;
            32'hB0001DAC: data = 32'd107;
            32'hB0001DB0: data = 32'd108;
            32'hB0001DB4: data = 32'd109;
            32'hB0001DB8: data = 32'd110;
            32'hB0001DBC: data = 32'd111;
            32'hB0001DC0: data = 32'd112;
            32'hB0001DC4: data = 32'd113;
            32'hB0001DC8: data = 32'd114;
            32'hB0001DCC: data = 32'd115;
            32'hB0001DD0: data = 32'd116;
            32'hB0001DD4: data = 32'd117;
            32'hB0001DD8: data = 32'd118;
            32'hB0001DDC: data = 32'd119;
            32'hB0001DE0: data = 32'd120;
            32'hB0001DE4: data = 32'd121;
            32'hB0001DE8: data = 32'd122;
            32'hB0001DEC: data = 32'd123;
            32'hB0001DF0: data = 32'd124;
            32'hB0001DF4: data = 32'd125;
            32'hB0001DF8: data = 32'd126;
            32'hB0001DFC: data = 32'd127;
            32'hB0001E00: data = 32'd128;
            32'hB0001E04: data = 32'd129;
            32'hB0001E08: data = 32'd130;
            32'hB0001E0C: data = 32'd131;
            32'hB0001E10: data = 32'd132;
            32'hB0001E14: data = 32'd133;
            32'hB0001E18: data = 32'd134;
            32'hB0001E1C: data = 32'd135;
            32'hB0001E20: data = 32'd136;
            32'hB0001E24: data = 32'd137;
            32'hB0001E28: data = 32'd138;
            32'hB0001E2C: data = 32'd139;
            32'hB0001E30: data = 32'd140;
            32'hB0001E34: data = 32'd141;
            32'hB0001E38: data = 32'd142;
            32'hB0001E3C: data = 32'd143;
            32'hB0001E40: data = 32'd144;
            32'hB0001E44: data = 32'd145;
            32'hB0001E48: data = 32'd146;
            32'hB0001E4C: data = 32'd147;
            32'hB0001E50: data = 32'd148;
            32'hB0001E54: data = 32'd149;
            32'hB0001E58: data = 32'd150;
            32'hB0001E5C: data = 32'd151;
            32'hB0001E60: data = 32'd152;
            32'hB0001E64: data = 32'd153;
            32'hB0001E68: data = 32'd154;
            32'hB0001E6C: data = 32'd155;
            32'hB0001E70: data = 32'd156;
            32'hB0001E74: data = 32'd157;
            32'hB0001E78: data = 32'd158;
            32'hB0001E7C: data = 32'd159;
            32'hB0001E80: data = 32'd160;
            32'hB0001E84: data = 32'd161;
            32'hB0001E88: data = 32'd162;
            32'hB0001E8C: data = 32'd163;
            32'hB0001E90: data = 32'd164;
            32'hB0001E94: data = 32'd165;
            32'hB0001E98: data = 32'd166;
            32'hB0001E9C: data = 32'd167;
            32'hB0001EA0: data = 32'd168;
            32'hB0001EA4: data = 32'd169;
            32'hB0001EA8: data = 32'd170;
            32'hB0001EAC: data = 32'd171;
            32'hB0001EB0: data = 32'd172;
            32'hB0001EB4: data = 32'd173;
            32'hB0001EB8: data = 32'd174;
            32'hB0001EBC: data = 32'd175;
            32'hB0001EC0: data = 32'd176;
            32'hB0001EC4: data = 32'd177;
            32'hB0001EC8: data = 32'd178;
            32'hB0001ECC: data = 32'd179;
            32'hB0001ED0: data = 32'd180;
            32'hB0001ED4: data = 32'd181;
            32'hB0001ED8: data = 32'd182;
            32'hB0001EDC: data = 32'd183;
            32'hB0001EE0: data = 32'd184;
            32'hB0001EE4: data = 32'd185;
            32'hB0001EE8: data = 32'd186;
            32'hB0001EEC: data = 32'd187;
            32'hB0001EF0: data = 32'd188;
            32'hB0001EF4: data = 32'd189;
            32'hB0001EF8: data = 32'd190;
            32'hB0001EFC: data = 32'd191;
            32'hB0001F00: data = 32'd192;
            32'hB0001F04: data = 32'd193;
            32'hB0001F08: data = 32'd194;
            32'hB0001F0C: data = 32'd195;
            32'hB0001F10: data = 32'd196;
            32'hB0001F14: data = 32'd197;
            32'hB0001F18: data = 32'd198;
            32'hB0001F1C: data = 32'd199;
            32'hB0001F20: data = 32'd200;
            32'hB0001F24: data = 32'd201;
            32'hB0001F28: data = 32'd202;
            32'hB0001F2C: data = 32'd203;
            32'hB0001F30: data = 32'd204;
            32'hB0001F34: data = 32'd205;
            32'hB0001F38: data = 32'd206;
            32'hB0001F3C: data = 32'd207;
            default: data = 32'd0;
        endcase
    end

endmodule

