module LUT_neg15degrees (
    input logic [9:0] counter,        // Counter ranging from 0 to 783
    output logic [11:0] address_offset       // Rotated address output
);

    always_comb begin
      case (counter) 
        

        10'b 0000000000 :   address_offset = 12'b 000000000000 ;
        10'b 0000000001 :   address_offset = 12'b 000000000000 ;
        10'b 0000000010 :   address_offset = 12'b 000000000000 ;
        10'b 0000000011 :   address_offset = 12'b 000101010000 ;
        10'b 0000000100 :   address_offset = 12'b 000101010100 ;
        10'b 0000000101 :   address_offset = 12'b 000101011000 ;
        10'b 0000000110 :   address_offset = 12'b 000101011100 ;
        10'b 0000000111 :   address_offset = 12'b 000011110000 ;
        10'b 0000001000 :   address_offset = 12'b 000011110100 ;
        10'b 0000001001 :   address_offset = 12'b 000011111000 ;
        10'b 0000001010 :   address_offset = 12'b 000011111100 ;
        10'b 0000001011 :   address_offset = 12'b 000010001100 ;
        10'b 0000001100 :   address_offset = 12'b 000010010000 ;
        10'b 0000001101 :   address_offset = 12'b 000010010100 ;
        10'b 0000001110 :   address_offset = 12'b 000000101000 ;
        10'b 0000001111 :   address_offset = 12'b 000000101100 ;
        10'b 0000010000 :   address_offset = 12'b 000000110000 ;
        10'b 0000010001 :   address_offset = 12'b 000000110100 ;
        10'b 0000010010 :   address_offset = 12'b 000000000000 ;
        10'b 0000010011 :   address_offset = 12'b 000000000000 ;
        10'b 0000010100 :   address_offset = 12'b 000000000000 ;
        10'b 0000010101 :   address_offset = 12'b 000000000000 ;
        10'b 0000010110 :   address_offset = 12'b 000000000000 ;
        10'b 0000010111 :   address_offset = 12'b 000000000000 ;
        10'b 0000011000 :   address_offset = 12'b 000000000000 ;
        10'b 0000011001 :   address_offset = 12'b 000000000000 ;
        10'b 0000011010 :   address_offset = 12'b 000000000000 ;
        10'b 0000011011 :   address_offset = 12'b 000000000000 ;
        10'b 0000011100 :   address_offset = 12'b 000000000000 ;
        10'b 0000011101 :   address_offset = 12'b 000000000000 ;
        10'b 0000011110 :   address_offset = 12'b 000000000000 ;
        10'b 0000011111 :   address_offset = 12'b 000111000000 ;
        10'b 0000100000 :   address_offset = 12'b 000111000100 ;
        10'b 0000100001 :   address_offset = 12'b 000111001000 ;
        10'b 0000100010 :   address_offset = 12'b 000111001100 ;
        10'b 0000100011 :   address_offset = 12'b 000101100000 ;
        10'b 0000100100 :   address_offset = 12'b 000101100100 ;
        10'b 0000100101 :   address_offset = 12'b 000101101000 ;
        10'b 0000100110 :   address_offset = 12'b 000011111100 ;
        10'b 0000100111 :   address_offset = 12'b 000100000000 ;
        10'b 0000101000 :   address_offset = 12'b 000100000100 ;
        10'b 0000101001 :   address_offset = 12'b 000100001000 ;
        10'b 0000101010 :   address_offset = 12'b 000010011100 ;
        10'b 0000101011 :   address_offset = 12'b 000010100000 ;
        10'b 0000101100 :   address_offset = 12'b 000010100100 ;
        10'b 0000101101 :   address_offset = 12'b 000010101000 ;
        10'b 0000101110 :   address_offset = 12'b 000000111000 ;
        10'b 0000101111 :   address_offset = 12'b 000000111100 ;
        10'b 0000110000 :   address_offset = 12'b 000001000000 ;
        10'b 0000110001 :   address_offset = 12'b 000001000100 ;
        10'b 0000110010 :   address_offset = 12'b 000000000000 ;
        10'b 0000110011 :   address_offset = 12'b 000000000000 ;
        10'b 0000110100 :   address_offset = 12'b 000000000000 ;
        10'b 0000110101 :   address_offset = 12'b 000000000000 ;
        10'b 0000110110 :   address_offset = 12'b 000000000000 ;
        10'b 0000110111 :   address_offset = 12'b 000000000000 ;
        10'b 0000111000 :   address_offset = 12'b 000000000000 ;
        10'b 0000111001 :   address_offset = 12'b 000000000000 ;
        10'b 0000111010 :   address_offset = 12'b 000000000000 ;
        10'b 0000111011 :   address_offset = 12'b 001000110000 ;
        10'b 0000111100 :   address_offset = 12'b 001000110100 ;
        10'b 0000111101 :   address_offset = 12'b 001000111000 ;
        10'b 0000111110 :   address_offset = 12'b 000111001100 ;
        10'b 0000111111 :   address_offset = 12'b 000111010000 ;
        10'b 0001000000 :   address_offset = 12'b 000111010100 ;
        10'b 0001000001 :   address_offset = 12'b 000111011000 ;
        10'b 0001000010 :   address_offset = 12'b 000101101100 ;
        10'b 0001000011 :   address_offset = 12'b 000101110000 ;
        10'b 0001000100 :   address_offset = 12'b 000101110100 ;
        10'b 0001000101 :   address_offset = 12'b 000101111000 ;
        10'b 0001000110 :   address_offset = 12'b 000100001100 ;
        10'b 0001000111 :   address_offset = 12'b 000100010000 ;
        10'b 0001001000 :   address_offset = 12'b 000100010100 ;
        10'b 0001001001 :   address_offset = 12'b 000100011000 ;
        10'b 0001001010 :   address_offset = 12'b 000010101100 ;
        10'b 0001001011 :   address_offset = 12'b 000010110000 ;
        10'b 0001001100 :   address_offset = 12'b 000010110100 ;
        10'b 0001001101 :   address_offset = 12'b 000010111000 ;
        10'b 0001001110 :   address_offset = 12'b 000001001100 ;
        10'b 0001001111 :   address_offset = 12'b 000001010000 ;
        10'b 0001010000 :   address_offset = 12'b 000001010100 ;
        10'b 0001010001 :   address_offset = 12'b 000001011000 ;
        10'b 0001010010 :   address_offset = 12'b 000000000000 ;
        10'b 0001010011 :   address_offset = 12'b 000000000000 ;
        10'b 0001010100 :   address_offset = 12'b 000000000000 ;
        10'b 0001010101 :   address_offset = 12'b 000000000000 ;
        10'b 0001010110 :   address_offset = 12'b 001010100000 ;
        10'b 0001010111 :   address_offset = 12'b 001010100100 ;
        10'b 0001011000 :   address_offset = 12'b 001010100100 ;
        10'b 0001011001 :   address_offset = 12'b 001010101000 ;
        10'b 0001011010 :   address_offset = 12'b 001000111100 ;
        10'b 0001011011 :   address_offset = 12'b 001001000000 ;
        10'b 0001011100 :   address_offset = 12'b 001001000100 ;
        10'b 0001011101 :   address_offset = 12'b 001001001000 ;
        10'b 0001011110 :   address_offset = 12'b 000111011100 ;
        10'b 0001011111 :   address_offset = 12'b 000111100000 ;
        10'b 0001100000 :   address_offset = 12'b 000111100100 ;
        10'b 0001100001 :   address_offset = 12'b 000111101000 ;
        10'b 0001100010 :   address_offset = 12'b 000101111100 ;
        10'b 0001100011 :   address_offset = 12'b 000110000000 ;
        10'b 0001100100 :   address_offset = 12'b 000110000100 ;
        10'b 0001100101 :   address_offset = 12'b 000110001000 ;
        10'b 0001100110 :   address_offset = 12'b 000100011100 ;
        10'b 0001100111 :   address_offset = 12'b 000100100000 ;
        10'b 0001101000 :   address_offset = 12'b 000100100100 ;
        10'b 0001101001 :   address_offset = 12'b 000100101000 ;
        10'b 0001101010 :   address_offset = 12'b 000010111100 ;
        10'b 0001101011 :   address_offset = 12'b 000011000000 ;
        10'b 0001101100 :   address_offset = 12'b 000011000100 ;
        10'b 0001101101 :   address_offset = 12'b 000011001000 ;
        10'b 0001101110 :   address_offset = 12'b 000001011100 ;
        10'b 0001101111 :   address_offset = 12'b 000001100000 ;
        10'b 0001110000 :   address_offset = 12'b 000000000000 ;
        10'b 0001110001 :   address_offset = 12'b 000000000000 ;
        10'b 0001110010 :   address_offset = 12'b 001100010000 ;
        10'b 0001110011 :   address_offset = 12'b 001100010100 ;
        10'b 0001110100 :   address_offset = 12'b 001100011000 ;
        10'b 0001110101 :   address_offset = 12'b 001100011100 ;
        10'b 0001110110 :   address_offset = 12'b 001010110000 ;
        10'b 0001110111 :   address_offset = 12'b 001010110100 ;
        10'b 0001111000 :   address_offset = 12'b 001010111000 ;
        10'b 0001111001 :   address_offset = 12'b 001010111100 ;
        10'b 0001111010 :   address_offset = 12'b 001001010000 ;
        10'b 0001111011 :   address_offset = 12'b 001001010100 ;
        10'b 0001111100 :   address_offset = 12'b 001001010100 ;
        10'b 0001111101 :   address_offset = 12'b 001001011000 ;
        10'b 0001111110 :   address_offset = 12'b 000111101100 ;
        10'b 0001111111 :   address_offset = 12'b 000111110000 ;
        10'b 0010000000 :   address_offset = 12'b 000111110100 ;
        10'b 0010000001 :   address_offset = 12'b 000111111000 ;
        10'b 0010000010 :   address_offset = 12'b 000110001100 ;
        10'b 0010000011 :   address_offset = 12'b 000110010000 ;
        10'b 0010000100 :   address_offset = 12'b 000110010100 ;
        10'b 0010000101 :   address_offset = 12'b 000110011000 ;
        10'b 0010000110 :   address_offset = 12'b 000100101100 ;
        10'b 0010000111 :   address_offset = 12'b 000100110000 ;
        10'b 0010001000 :   address_offset = 12'b 000100110100 ;
        10'b 0010001001 :   address_offset = 12'b 000011001000 ;
        10'b 0010001010 :   address_offset = 12'b 000011001100 ;
        10'b 0010001011 :   address_offset = 12'b 000011010000 ;
        10'b 0010001100 :   address_offset = 12'b 000000000000 ;
        10'b 0010001101 :   address_offset = 12'b 000000000000 ;
        10'b 0010001110 :   address_offset = 12'b 001110000000 ;
        10'b 0010001111 :   address_offset = 12'b 001110000100 ;
        10'b 0010010000 :   address_offset = 12'b 001110001000 ;
        10'b 0010010001 :   address_offset = 12'b 001110001100 ;
        10'b 0010010010 :   address_offset = 12'b 001100100000 ;
        10'b 0010010011 :   address_offset = 12'b 001100100100 ;
        10'b 0010010100 :   address_offset = 12'b 001100101000 ;
        10'b 0010010101 :   address_offset = 12'b 001100101100 ;
        10'b 0010010110 :   address_offset = 12'b 001011000000 ;
        10'b 0010010111 :   address_offset = 12'b 001011000100 ;
        10'b 0010011000 :   address_offset = 12'b 001011001000 ;
        10'b 0010011001 :   address_offset = 12'b 001011001100 ;
        10'b 0010011010 :   address_offset = 12'b 001001100000 ;
        10'b 0010011011 :   address_offset = 12'b 001001100100 ;
        10'b 0010011100 :   address_offset = 12'b 001001101000 ;
        10'b 0010011101 :   address_offset = 12'b 001001101100 ;
        10'b 0010011110 :   address_offset = 12'b 001000000000 ;
        10'b 0010011111 :   address_offset = 12'b 001000000100 ;
        10'b 0010100000 :   address_offset = 12'b 001000000100 ;
        10'b 0010100001 :   address_offset = 12'b 000110011000 ;
        10'b 0010100010 :   address_offset = 12'b 000110011100 ;
        10'b 0010100011 :   address_offset = 12'b 000110100000 ;
        10'b 0010100100 :   address_offset = 12'b 000110100100 ;
        10'b 0010100101 :   address_offset = 12'b 000100111000 ;
        10'b 0010100110 :   address_offset = 12'b 000100111100 ;
        10'b 0010100111 :   address_offset = 12'b 000101000000 ;
        10'b 0010101000 :   address_offset = 12'b 000000000000 ;
        10'b 0010101001 :   address_offset = 12'b 000000000000 ;
        10'b 0010101010 :   address_offset = 12'b 001111110000 ;
        10'b 0010101011 :   address_offset = 12'b 001111110100 ;
        10'b 0010101100 :   address_offset = 12'b 001111111000 ;
        10'b 0010101101 :   address_offset = 12'b 001111111100 ;
        10'b 0010101110 :   address_offset = 12'b 001110010000 ;
        10'b 0010101111 :   address_offset = 12'b 001110010100 ;
        10'b 0010110000 :   address_offset = 12'b 001110011000 ;
        10'b 0010110001 :   address_offset = 12'b 001110011100 ;
        10'b 0010110010 :   address_offset = 12'b 001100110000 ;
        10'b 0010110011 :   address_offset = 12'b 001100110100 ;
        10'b 0010110100 :   address_offset = 12'b 001100111000 ;
        10'b 0010110101 :   address_offset = 12'b 001100111100 ;
        10'b 0010110110 :   address_offset = 12'b 001011010000 ;
        10'b 0010110111 :   address_offset = 12'b 001011010100 ;
        10'b 0010111000 :   address_offset = 12'b 001011011000 ;
        10'b 0010111001 :   address_offset = 12'b 001001101100 ;
        10'b 0010111010 :   address_offset = 12'b 001001110000 ;
        10'b 0010111011 :   address_offset = 12'b 001001110100 ;
        10'b 0010111100 :   address_offset = 12'b 001001111000 ;
        10'b 0010111101 :   address_offset = 12'b 001000001100 ;
        10'b 0010111110 :   address_offset = 12'b 001000010000 ;
        10'b 0010111111 :   address_offset = 12'b 001000010100 ;
        10'b 0011000000 :   address_offset = 12'b 001000011000 ;
        10'b 0011000001 :   address_offset = 12'b 000110101100 ;
        10'b 0011000010 :   address_offset = 12'b 000110110000 ;
        10'b 0011000011 :   address_offset = 12'b 000110110000 ;
        10'b 0011000100 :   address_offset = 12'b 000000000000 ;
        10'b 0011000101 :   address_offset = 12'b 010011010000 ;
        10'b 0011000110 :   address_offset = 12'b 010001100100 ;
        10'b 0011000111 :   address_offset = 12'b 010001101000 ;
        10'b 0011001000 :   address_offset = 12'b 010001101100 ;
        10'b 0011001001 :   address_offset = 12'b 010001101100 ;
        10'b 0011001010 :   address_offset = 12'b 010000000000 ;
        10'b 0011001011 :   address_offset = 12'b 010000000100 ;
        10'b 0011001100 :   address_offset = 12'b 010000001000 ;
        10'b 0011001101 :   address_offset = 12'b 010000001100 ;
        10'b 0011001110 :   address_offset = 12'b 001110100000 ;
        10'b 0011001111 :   address_offset = 12'b 001110100100 ;
        10'b 0011010000 :   address_offset = 12'b 001110101000 ;
        10'b 0011010001 :   address_offset = 12'b 001100111100 ;
        10'b 0011010010 :   address_offset = 12'b 001101000000 ;
        10'b 0011010011 :   address_offset = 12'b 001101000100 ;
        10'b 0011010100 :   address_offset = 12'b 001101001000 ;
        10'b 0011010101 :   address_offset = 12'b 001011011100 ;
        10'b 0011010110 :   address_offset = 12'b 001011100000 ;
        10'b 0011010111 :   address_offset = 12'b 001011100100 ;
        10'b 0011011000 :   address_offset = 12'b 001011101000 ;
        10'b 0011011001 :   address_offset = 12'b 001001111100 ;
        10'b 0011011010 :   address_offset = 12'b 001010000000 ;
        10'b 0011011011 :   address_offset = 12'b 001010000100 ;
        10'b 0011011100 :   address_offset = 12'b 001010001000 ;
        10'b 0011011101 :   address_offset = 12'b 001000011100 ;
        10'b 0011011110 :   address_offset = 12'b 001000100000 ;
        10'b 0011011111 :   address_offset = 12'b 001000100100 ;
        10'b 0011100000 :   address_offset = 12'b 000000000000 ;
        10'b 0011100001 :   address_offset = 12'b 010101000000 ;
        10'b 0011100010 :   address_offset = 12'b 010011010100 ;
        10'b 0011100011 :   address_offset = 12'b 010011011000 ;
        10'b 0011100100 :   address_offset = 12'b 010011011100 ;
        10'b 0011100101 :   address_offset = 12'b 010011100000 ;
        10'b 0011100110 :   address_offset = 12'b 010001110100 ;
        10'b 0011100111 :   address_offset = 12'b 010001111000 ;
        10'b 0011101000 :   address_offset = 12'b 010001111100 ;
        10'b 0011101001 :   address_offset = 12'b 010000010000 ;
        10'b 0011101010 :   address_offset = 12'b 010000010100 ;
        10'b 0011101011 :   address_offset = 12'b 010000011000 ;
        10'b 0011101100 :   address_offset = 12'b 010000011100 ;
        10'b 0011101101 :   address_offset = 12'b 001110101100 ;
        10'b 0011101110 :   address_offset = 12'b 001110110000 ;
        10'b 0011101111 :   address_offset = 12'b 001110110100 ;
        10'b 0011110000 :   address_offset = 12'b 001110111000 ;
        10'b 0011110001 :   address_offset = 12'b 001101001100 ;
        10'b 0011110010 :   address_offset = 12'b 001101010000 ;
        10'b 0011110011 :   address_offset = 12'b 001101010100 ;
        10'b 0011110100 :   address_offset = 12'b 001101011000 ;
        10'b 0011110101 :   address_offset = 12'b 001011101100 ;
        10'b 0011110110 :   address_offset = 12'b 001011110000 ;
        10'b 0011110111 :   address_offset = 12'b 001011110100 ;
        10'b 0011111000 :   address_offset = 12'b 001011111000 ;
        10'b 0011111001 :   address_offset = 12'b 001010001100 ;
        10'b 0011111010 :   address_offset = 12'b 001010010000 ;
        10'b 0011111011 :   address_offset = 12'b 001010010100 ;
        10'b 0011111100 :   address_offset = 12'b 000000000000 ;
        10'b 0011111101 :   address_offset = 12'b 010110110000 ;
        10'b 0011111110 :   address_offset = 12'b 010101000100 ;
        10'b 0011111111 :   address_offset = 12'b 010101001000 ;
        10'b 0100000000 :   address_offset = 12'b 010101001100 ;
        10'b 0100000001 :   address_offset = 12'b 010011100000 ;
        10'b 0100000010 :   address_offset = 12'b 010011100100 ;
        10'b 0100000011 :   address_offset = 12'b 010011101000 ;
        10'b 0100000100 :   address_offset = 12'b 010011101100 ;
        10'b 0100000101 :   address_offset = 12'b 010010000000 ;
        10'b 0100000110 :   address_offset = 12'b 010010000100 ;
        10'b 0100000111 :   address_offset = 12'b 010010001000 ;
        10'b 0100001000 :   address_offset = 12'b 010010001100 ;
        10'b 0100001001 :   address_offset = 12'b 010000100000 ;
        10'b 0100001010 :   address_offset = 12'b 010000100100 ;
        10'b 0100001011 :   address_offset = 12'b 010000101000 ;
        10'b 0100001100 :   address_offset = 12'b 010000101100 ;
        10'b 0100001101 :   address_offset = 12'b 001111000000 ;
        10'b 0100001110 :   address_offset = 12'b 001111000100 ;
        10'b 0100001111 :   address_offset = 12'b 001111001000 ;
        10'b 0100010000 :   address_offset = 12'b 001111001100 ;
        10'b 0100010001 :   address_offset = 12'b 001101011100 ;
        10'b 0100010010 :   address_offset = 12'b 001101100000 ;
        10'b 0100010011 :   address_offset = 12'b 001101100100 ;
        10'b 0100010100 :   address_offset = 12'b 001101101000 ;
        10'b 0100010101 :   address_offset = 12'b 001011111100 ;
        10'b 0100010110 :   address_offset = 12'b 001100000000 ;
        10'b 0100010111 :   address_offset = 12'b 001100000100 ;
        10'b 0100011000 :   address_offset = 12'b 000000000000 ;
        10'b 0100011001 :   address_offset = 12'b 011000100000 ;
        10'b 0100011010 :   address_offset = 12'b 010110110100 ;
        10'b 0100011011 :   address_offset = 12'b 010110111000 ;
        10'b 0100011100 :   address_offset = 12'b 010110111100 ;
        10'b 0100011101 :   address_offset = 12'b 010101010000 ;
        10'b 0100011110 :   address_offset = 12'b 010101010100 ;
        10'b 0100011111 :   address_offset = 12'b 010101011000 ;
        10'b 0100100000 :   address_offset = 12'b 010101011100 ;
        10'b 0100100001 :   address_offset = 12'b 010011110000 ;
        10'b 0100100010 :   address_offset = 12'b 010011110100 ;
        10'b 0100100011 :   address_offset = 12'b 010011111000 ;
        10'b 0100100100 :   address_offset = 12'b 010011111100 ;
        10'b 0100100101 :   address_offset = 12'b 010010010000 ;
        10'b 0100100110 :   address_offset = 12'b 010010010100 ;
        10'b 0100100111 :   address_offset = 12'b 010010011000 ;
        10'b 0100101000 :   address_offset = 12'b 010010011100 ;
        10'b 0100101001 :   address_offset = 12'b 010000110000 ;
        10'b 0100101010 :   address_offset = 12'b 010000110100 ;
        10'b 0100101011 :   address_offset = 12'b 010000111000 ;
        10'b 0100101100 :   address_offset = 12'b 010000111100 ;
        10'b 0100101101 :   address_offset = 12'b 001111010000 ;
        10'b 0100101110 :   address_offset = 12'b 001111010100 ;
        10'b 0100101111 :   address_offset = 12'b 001111011000 ;
        10'b 0100110000 :   address_offset = 12'b 001111011100 ;
        10'b 0100110001 :   address_offset = 12'b 001101110000 ;
        10'b 0100110010 :   address_offset = 12'b 001101110100 ;
        10'b 0100110011 :   address_offset = 12'b 001101111000 ;
        10'b 0100110100 :   address_offset = 12'b 011010010000 ;
        10'b 0100110101 :   address_offset = 12'b 011000100100 ;
        10'b 0100110110 :   address_offset = 12'b 011000101000 ;
        10'b 0100110111 :   address_offset = 12'b 011000101100 ;
        10'b 0100111000 :   address_offset = 12'b 011000110000 ;
        10'b 0100111001 :   address_offset = 12'b 010111000100 ;
        10'b 0100111010 :   address_offset = 12'b 010111000100 ;
        10'b 0100111011 :   address_offset = 12'b 010111001000 ;
        10'b 0100111100 :   address_offset = 12'b 010111001100 ;
        10'b 0100111101 :   address_offset = 12'b 010101100000 ;
        10'b 0100111110 :   address_offset = 12'b 010101100100 ;
        10'b 0100111111 :   address_offset = 12'b 010101101000 ;
        10'b 0101000000 :   address_offset = 12'b 010101101100 ;
        10'b 0101000001 :   address_offset = 12'b 010100000000 ;
        10'b 0101000010 :   address_offset = 12'b 010100000100 ;
        10'b 0101000011 :   address_offset = 12'b 010100001000 ;
        10'b 0101000100 :   address_offset = 12'b 010100001100 ;
        10'b 0101000101 :   address_offset = 12'b 010010100000 ;
        10'b 0101000110 :   address_offset = 12'b 010010100100 ;
        10'b 0101000111 :   address_offset = 12'b 010010101000 ;
        10'b 0101001000 :   address_offset = 12'b 010010101100 ;
        10'b 0101001001 :   address_offset = 12'b 010001000000 ;
        10'b 0101001010 :   address_offset = 12'b 010001000100 ;
        10'b 0101001011 :   address_offset = 12'b 010001001000 ;
        10'b 0101001100 :   address_offset = 12'b 010001001100 ;
        10'b 0101001101 :   address_offset = 12'b 001111100000 ;
        10'b 0101001110 :   address_offset = 12'b 001111100100 ;
        10'b 0101001111 :   address_offset = 12'b 001111101000 ;
        10'b 0101010000 :   address_offset = 12'b 011100000000 ;
        10'b 0101010001 :   address_offset = 12'b 011010010100 ;
        10'b 0101010010 :   address_offset = 12'b 011010011000 ;
        10'b 0101010011 :   address_offset = 12'b 011010011100 ;
        10'b 0101010100 :   address_offset = 12'b 011010100000 ;
        10'b 0101010101 :   address_offset = 12'b 011000110100 ;
        10'b 0101010110 :   address_offset = 12'b 011000111000 ;
        10'b 0101010111 :   address_offset = 12'b 011000111100 ;
        10'b 0101011000 :   address_offset = 12'b 011001000000 ;
        10'b 0101011001 :   address_offset = 12'b 010111010100 ;
        10'b 0101011010 :   address_offset = 12'b 010111011000 ;
        10'b 0101011011 :   address_offset = 12'b 010111011100 ;
        10'b 0101011100 :   address_offset = 12'b 010111100000 ;
        10'b 0101011101 :   address_offset = 12'b 010101110100 ;
        10'b 0101011110 :   address_offset = 12'b 010101110100 ;
        10'b 0101011111 :   address_offset = 12'b 010101111000 ;
        10'b 0101100000 :   address_offset = 12'b 010101111100 ;
        10'b 0101100001 :   address_offset = 12'b 010100010000 ;
        10'b 0101100010 :   address_offset = 12'b 010100010100 ;
        10'b 0101100011 :   address_offset = 12'b 010100011000 ;
        10'b 0101100100 :   address_offset = 12'b 010100011100 ;
        10'b 0101100101 :   address_offset = 12'b 010010110000 ;
        10'b 0101100110 :   address_offset = 12'b 010010110100 ;
        10'b 0101100111 :   address_offset = 12'b 010010111000 ;
        10'b 0101101000 :   address_offset = 12'b 010001001100 ;
        10'b 0101101001 :   address_offset = 12'b 010001010000 ;
        10'b 0101101010 :   address_offset = 12'b 010001010100 ;
        10'b 0101101011 :   address_offset = 12'b 010001011000 ;
        10'b 0101101100 :   address_offset = 12'b 011101110000 ;
        10'b 0101101101 :   address_offset = 12'b 011100000100 ;
        10'b 0101101110 :   address_offset = 12'b 011100001000 ;
        10'b 0101101111 :   address_offset = 12'b 011100001100 ;
        10'b 0101110000 :   address_offset = 12'b 011100010000 ;
        10'b 0101110001 :   address_offset = 12'b 011010100100 ;
        10'b 0101110010 :   address_offset = 12'b 011010101000 ;
        10'b 0101110011 :   address_offset = 12'b 011010101100 ;
        10'b 0101110100 :   address_offset = 12'b 011010110000 ;
        10'b 0101110101 :   address_offset = 12'b 011001000100 ;
        10'b 0101110110 :   address_offset = 12'b 011001001000 ;
        10'b 0101110111 :   address_offset = 12'b 011001001100 ;
        10'b 0101111000 :   address_offset = 12'b 011001010000 ;
        10'b 0101111001 :   address_offset = 12'b 010111100100 ;
        10'b 0101111010 :   address_offset = 12'b 010111101000 ;
        10'b 0101111011 :   address_offset = 12'b 010111101100 ;
        10'b 0101111100 :   address_offset = 12'b 010111110000 ;
        10'b 0101111101 :   address_offset = 12'b 010110000100 ;
        10'b 0101111110 :   address_offset = 12'b 010110001000 ;
        10'b 0101111111 :   address_offset = 12'b 010110001100 ;
        10'b 0110000000 :   address_offset = 12'b 010100100000 ;
        10'b 0110000001 :   address_offset = 12'b 010100100100 ;
        10'b 0110000010 :   address_offset = 12'b 010100100100 ;
        10'b 0110000011 :   address_offset = 12'b 010100101000 ;
        10'b 0110000100 :   address_offset = 12'b 010010111100 ;
        10'b 0110000101 :   address_offset = 12'b 010011000000 ;
        10'b 0110000110 :   address_offset = 12'b 010011000100 ;
        10'b 0110000111 :   address_offset = 12'b 010011001000 ;
        10'b 0110001000 :   address_offset = 12'b 011111100000 ;
        10'b 0110001001 :   address_offset = 12'b 011101110100 ;
        10'b 0110001010 :   address_offset = 12'b 011101111000 ;
        10'b 0110001011 :   address_offset = 12'b 011101111100 ;
        10'b 0110001100 :   address_offset = 12'b 011110000000 ;
        10'b 0110001101 :   address_offset = 12'b 011100010100 ;
        10'b 0110001110 :   address_offset = 12'b 011100011000 ;
        10'b 0110001111 :   address_offset = 12'b 011100011100 ;
        10'b 0110010000 :   address_offset = 12'b 011100100000 ;
        10'b 0110010001 :   address_offset = 12'b 011010110100 ;
        10'b 0110010010 :   address_offset = 12'b 011010111000 ;
        10'b 0110010011 :   address_offset = 12'b 011010111100 ;
        10'b 0110010100 :   address_offset = 12'b 011011000000 ;
        10'b 0110010101 :   address_offset = 12'b 011001010100 ;
        10'b 0110010110 :   address_offset = 12'b 011001011000 ;
        10'b 0110010111 :   address_offset = 12'b 011001011100 ;
        10'b 0110011000 :   address_offset = 12'b 010111110000 ;
        10'b 0110011001 :   address_offset = 12'b 010111110100 ;
        10'b 0110011010 :   address_offset = 12'b 010111111000 ;
        10'b 0110011011 :   address_offset = 12'b 010111111100 ;
        10'b 0110011100 :   address_offset = 12'b 010110010000 ;
        10'b 0110011101 :   address_offset = 12'b 010110010100 ;
        10'b 0110011110 :   address_offset = 12'b 010110011000 ;
        10'b 0110011111 :   address_offset = 12'b 010110011100 ;
        10'b 0110100000 :   address_offset = 12'b 010100110000 ;
        10'b 0110100001 :   address_offset = 12'b 010100110100 ;
        10'b 0110100010 :   address_offset = 12'b 010100111000 ;
        10'b 0110100011 :   address_offset = 12'b 010100111100 ;
        10'b 0110100100 :   address_offset = 12'b 100001010100 ;
        10'b 0110100101 :   address_offset = 12'b 011111101000 ;
        10'b 0110100110 :   address_offset = 12'b 011111101100 ;
        10'b 0110100111 :   address_offset = 12'b 011111110000 ;
        10'b 0110101000 :   address_offset = 12'b 011111110100 ;
        10'b 0110101001 :   address_offset = 12'b 011110001000 ;
        10'b 0110101010 :   address_offset = 12'b 011110001100 ;
        10'b 0110101011 :   address_offset = 12'b 011110001100 ;
        10'b 0110101100 :   address_offset = 12'b 011110010000 ;
        10'b 0110101101 :   address_offset = 12'b 011100100100 ;
        10'b 0110101110 :   address_offset = 12'b 011100101000 ;
        10'b 0110101111 :   address_offset = 12'b 011100101100 ;
        10'b 0110110000 :   address_offset = 12'b 011011000000 ;
        10'b 0110110001 :   address_offset = 12'b 011011000100 ;
        10'b 0110110010 :   address_offset = 12'b 011011001000 ;
        10'b 0110110011 :   address_offset = 12'b 011011001100 ;
        10'b 0110110100 :   address_offset = 12'b 011001100000 ;
        10'b 0110110101 :   address_offset = 12'b 011001100100 ;
        10'b 0110110110 :   address_offset = 12'b 011001101000 ;
        10'b 0110110111 :   address_offset = 12'b 011001101100 ;
        10'b 0110111000 :   address_offset = 12'b 011000000000 ;
        10'b 0110111001 :   address_offset = 12'b 011000000100 ;
        10'b 0110111010 :   address_offset = 12'b 011000001000 ;
        10'b 0110111011 :   address_offset = 12'b 011000001100 ;
        10'b 0110111100 :   address_offset = 12'b 010110100000 ;
        10'b 0110111101 :   address_offset = 12'b 010110100100 ;
        10'b 0110111110 :   address_offset = 12'b 010110101000 ;
        10'b 0110111111 :   address_offset = 12'b 010110101100 ;
        10'b 0111000000 :   address_offset = 12'b 100011000100 ;
        10'b 0111000001 :   address_offset = 12'b 100001011000 ;
        10'b 0111000010 :   address_offset = 12'b 100001011100 ;
        10'b 0111000011 :   address_offset = 12'b 100001100000 ;
        10'b 0111000100 :   address_offset = 12'b 100001100100 ;
        10'b 0111000101 :   address_offset = 12'b 011111111000 ;
        10'b 0111000110 :   address_offset = 12'b 011111111100 ;
        10'b 0111000111 :   address_offset = 12'b 100000000000 ;
        10'b 0111001000 :   address_offset = 12'b 011110010100 ;
        10'b 0111001001 :   address_offset = 12'b 011110011000 ;
        10'b 0111001010 :   address_offset = 12'b 011110011100 ;
        10'b 0111001011 :   address_offset = 12'b 011110100000 ;
        10'b 0111001100 :   address_offset = 12'b 011100110100 ;
        10'b 0111001101 :   address_offset = 12'b 011100111000 ;
        10'b 0111001110 :   address_offset = 12'b 011100111100 ;
        10'b 0111001111 :   address_offset = 12'b 011100111100 ;
        10'b 0111010000 :   address_offset = 12'b 011011010000 ;
        10'b 0111010001 :   address_offset = 12'b 011011010100 ;
        10'b 0111010010 :   address_offset = 12'b 011011011000 ;
        10'b 0111010011 :   address_offset = 12'b 011011011100 ;
        10'b 0111010100 :   address_offset = 12'b 011001110000 ;
        10'b 0111010101 :   address_offset = 12'b 011001110100 ;
        10'b 0111010110 :   address_offset = 12'b 011001111000 ;
        10'b 0111010111 :   address_offset = 12'b 011001111100 ;
        10'b 0111011000 :   address_offset = 12'b 011000010000 ;
        10'b 0111011001 :   address_offset = 12'b 011000010100 ;
        10'b 0111011010 :   address_offset = 12'b 011000011000 ;
        10'b 0111011011 :   address_offset = 12'b 011000011100 ;
        10'b 0111011100 :   address_offset = 12'b 100100110100 ;
        10'b 0111011101 :   address_offset = 12'b 100011001000 ;
        10'b 0111011110 :   address_offset = 12'b 100011001100 ;
        10'b 0111011111 :   address_offset = 12'b 100011010000 ;
        10'b 0111100000 :   address_offset = 12'b 100001100100 ;
        10'b 0111100001 :   address_offset = 12'b 100001101000 ;
        10'b 0111100010 :   address_offset = 12'b 100001101100 ;
        10'b 0111100011 :   address_offset = 12'b 100001110000 ;
        10'b 0111100100 :   address_offset = 12'b 100000000100 ;
        10'b 0111100101 :   address_offset = 12'b 100000001000 ;
        10'b 0111100110 :   address_offset = 12'b 100000001100 ;
        10'b 0111100111 :   address_offset = 12'b 100000010000 ;
        10'b 0111101000 :   address_offset = 12'b 011110100100 ;
        10'b 0111101001 :   address_offset = 12'b 011110101000 ;
        10'b 0111101010 :   address_offset = 12'b 011110101100 ;
        10'b 0111101011 :   address_offset = 12'b 011110110000 ;
        10'b 0111101100 :   address_offset = 12'b 011101000100 ;
        10'b 0111101101 :   address_offset = 12'b 011101001000 ;
        10'b 0111101110 :   address_offset = 12'b 011101001100 ;
        10'b 0111101111 :   address_offset = 12'b 011101010000 ;
        10'b 0111110000 :   address_offset = 12'b 011011100100 ;
        10'b 0111110001 :   address_offset = 12'b 011011101000 ;
        10'b 0111110010 :   address_offset = 12'b 011011101100 ;
        10'b 0111110011 :   address_offset = 12'b 011011101100 ;
        10'b 0111110100 :   address_offset = 12'b 011010000000 ;
        10'b 0111110101 :   address_offset = 12'b 011010000100 ;
        10'b 0111110110 :   address_offset = 12'b 011010001000 ;
        10'b 0111110111 :   address_offset = 12'b 011010001100 ;
        10'b 0111111000 :   address_offset = 12'b 100100111000 ;
        10'b 0111111001 :   address_offset = 12'b 100100111000 ;
        10'b 0111111010 :   address_offset = 12'b 100100111100 ;
        10'b 0111111011 :   address_offset = 12'b 100101000000 ;
        10'b 0111111100 :   address_offset = 12'b 100011010100 ;
        10'b 0111111101 :   address_offset = 12'b 100011011000 ;
        10'b 0111111110 :   address_offset = 12'b 100011011100 ;
        10'b 0111111111 :   address_offset = 12'b 100011100000 ;
        10'b 1000000000 :   address_offset = 12'b 100001110100 ;
        10'b 1000000001 :   address_offset = 12'b 100001111000 ;
        10'b 1000000010 :   address_offset = 12'b 100001111100 ;
        10'b 1000000011 :   address_offset = 12'b 100010000000 ;
        10'b 1000000100 :   address_offset = 12'b 100000010100 ;
        10'b 1000000101 :   address_offset = 12'b 100000011000 ;
        10'b 1000000110 :   address_offset = 12'b 100000011100 ;
        10'b 1000000111 :   address_offset = 12'b 100000100000 ;
        10'b 1000001000 :   address_offset = 12'b 011110110100 ;
        10'b 1000001001 :   address_offset = 12'b 011110111000 ;
        10'b 1000001010 :   address_offset = 12'b 011110111100 ;
        10'b 1000001011 :   address_offset = 12'b 011111000000 ;
        10'b 1000001100 :   address_offset = 12'b 011101010100 ;
        10'b 1000001101 :   address_offset = 12'b 011101011000 ;
        10'b 1000001110 :   address_offset = 12'b 011101011100 ;
        10'b 1000001111 :   address_offset = 12'b 011101100000 ;
        10'b 1000010000 :   address_offset = 12'b 011011110100 ;
        10'b 1000010001 :   address_offset = 12'b 011011111000 ;
        10'b 1000010010 :   address_offset = 12'b 011011111100 ;
        10'b 1000010011 :   address_offset = 12'b 000000000000 ;
        10'b 1000010100 :   address_offset = 12'b 100110101000 ;
        10'b 1000010101 :   address_offset = 12'b 100110101100 ;
        10'b 1000010110 :   address_offset = 12'b 100110110000 ;
        10'b 1000010111 :   address_offset = 12'b 100110110100 ;
        10'b 1000011000 :   address_offset = 12'b 100101001000 ;
        10'b 1000011001 :   address_offset = 12'b 100101001100 ;
        10'b 1000011010 :   address_offset = 12'b 100101010000 ;
        10'b 1000011011 :   address_offset = 12'b 100101010100 ;
        10'b 1000011100 :   address_offset = 12'b 100011100100 ;
        10'b 1000011101 :   address_offset = 12'b 100011101000 ;
        10'b 1000011110 :   address_offset = 12'b 100011101100 ;
        10'b 1000011111 :   address_offset = 12'b 100011110000 ;
        10'b 1000100000 :   address_offset = 12'b 100010000100 ;
        10'b 1000100001 :   address_offset = 12'b 100010001000 ;
        10'b 1000100010 :   address_offset = 12'b 100010001100 ;
        10'b 1000100011 :   address_offset = 12'b 100010010000 ;
        10'b 1000100100 :   address_offset = 12'b 100000100100 ;
        10'b 1000100101 :   address_offset = 12'b 100000101000 ;
        10'b 1000100110 :   address_offset = 12'b 100000101100 ;
        10'b 1000100111 :   address_offset = 12'b 100000110000 ;
        10'b 1000101000 :   address_offset = 12'b 011111000100 ;
        10'b 1000101001 :   address_offset = 12'b 011111001000 ;
        10'b 1000101010 :   address_offset = 12'b 011111001100 ;
        10'b 1000101011 :   address_offset = 12'b 011111010000 ;
        10'b 1000101100 :   address_offset = 12'b 011101100100 ;
        10'b 1000101101 :   address_offset = 12'b 011101101000 ;
        10'b 1000101110 :   address_offset = 12'b 011101101100 ;
        10'b 1000101111 :   address_offset = 12'b 000000000000 ;
        10'b 1000110000 :   address_offset = 12'b 101000011000 ;
        10'b 1000110001 :   address_offset = 12'b 101000011100 ;
        10'b 1000110010 :   address_offset = 12'b 101000100000 ;
        10'b 1000110011 :   address_offset = 12'b 101000100100 ;
        10'b 1000110100 :   address_offset = 12'b 100110111000 ;
        10'b 1000110101 :   address_offset = 12'b 100110111100 ;
        10'b 1000110110 :   address_offset = 12'b 100111000000 ;
        10'b 1000110111 :   address_offset = 12'b 100111000100 ;
        10'b 1000111000 :   address_offset = 12'b 100101011000 ;
        10'b 1000111001 :   address_offset = 12'b 100101011100 ;
        10'b 1000111010 :   address_offset = 12'b 100101100000 ;
        10'b 1000111011 :   address_offset = 12'b 100101100100 ;
        10'b 1000111100 :   address_offset = 12'b 100011111000 ;
        10'b 1000111101 :   address_offset = 12'b 100011111100 ;
        10'b 1000111110 :   address_offset = 12'b 100100000000 ;
        10'b 1000111111 :   address_offset = 12'b 100100000100 ;
        10'b 1001000000 :   address_offset = 12'b 100010010100 ;
        10'b 1001000001 :   address_offset = 12'b 100010011000 ;
        10'b 1001000010 :   address_offset = 12'b 100010011100 ;
        10'b 1001000011 :   address_offset = 12'b 100010100000 ;
        10'b 1001000100 :   address_offset = 12'b 100000110100 ;
        10'b 1001000101 :   address_offset = 12'b 100000111000 ;
        10'b 1001000110 :   address_offset = 12'b 100000111100 ;
        10'b 1001000111 :   address_offset = 12'b 011111010000 ;
        10'b 1001001000 :   address_offset = 12'b 011111010100 ;
        10'b 1001001001 :   address_offset = 12'b 011111011000 ;
        10'b 1001001010 :   address_offset = 12'b 011111011100 ;
        10'b 1001001011 :   address_offset = 12'b 000000000000 ;
        10'b 1001001100 :   address_offset = 12'b 101010001000 ;
        10'b 1001001101 :   address_offset = 12'b 101010001100 ;
        10'b 1001001110 :   address_offset = 12'b 101010010000 ;
        10'b 1001001111 :   address_offset = 12'b 101010010100 ;
        10'b 1001010000 :   address_offset = 12'b 101000101000 ;
        10'b 1001010001 :   address_offset = 12'b 101000101100 ;
        10'b 1001010010 :   address_offset = 12'b 101000110000 ;
        10'b 1001010011 :   address_offset = 12'b 101000110100 ;
        10'b 1001010100 :   address_offset = 12'b 100111001000 ;
        10'b 1001010101 :   address_offset = 12'b 100111001100 ;
        10'b 1001010110 :   address_offset = 12'b 100111010000 ;
        10'b 1001010111 :   address_offset = 12'b 100111010100 ;
        10'b 1001011000 :   address_offset = 12'b 100101101000 ;
        10'b 1001011001 :   address_offset = 12'b 100101101100 ;
        10'b 1001011010 :   address_offset = 12'b 100101110000 ;
        10'b 1001011011 :   address_offset = 12'b 100101110100 ;
        10'b 1001011100 :   address_offset = 12'b 100100001000 ;
        10'b 1001011101 :   address_offset = 12'b 100100001100 ;
        10'b 1001011110 :   address_offset = 12'b 100100010000 ;
        10'b 1001011111 :   address_offset = 12'b 100010100100 ;
        10'b 1001100000 :   address_offset = 12'b 100010101000 ;
        10'b 1001100001 :   address_offset = 12'b 100010101100 ;
        10'b 1001100010 :   address_offset = 12'b 100010110000 ;
        10'b 1001100011 :   address_offset = 12'b 100001000100 ;
        10'b 1001100100 :   address_offset = 12'b 100001000100 ;
        10'b 1001100101 :   address_offset = 12'b 100001001000 ;
        10'b 1001100110 :   address_offset = 12'b 100001001100 ;
        10'b 1001100111 :   address_offset = 12'b 000000000000 ;
        10'b 1001101000 :   address_offset = 12'b 101011111100 ;
        10'b 1001101001 :   address_offset = 12'b 101100000000 ;
        10'b 1001101010 :   address_offset = 12'b 101100000000 ;
        10'b 1001101011 :   address_offset = 12'b 101100000100 ;
        10'b 1001101100 :   address_offset = 12'b 101010011000 ;
        10'b 1001101101 :   address_offset = 12'b 101010011100 ;
        10'b 1001101110 :   address_offset = 12'b 101010100000 ;
        10'b 1001101111 :   address_offset = 12'b 101010100100 ;
        10'b 1001110000 :   address_offset = 12'b 101000111000 ;
        10'b 1001110001 :   address_offset = 12'b 101000111100 ;
        10'b 1001110010 :   address_offset = 12'b 101001000000 ;
        10'b 1001110011 :   address_offset = 12'b 101001000100 ;
        10'b 1001110100 :   address_offset = 12'b 100111011000 ;
        10'b 1001110101 :   address_offset = 12'b 100111011100 ;
        10'b 1001110110 :   address_offset = 12'b 100111100000 ;
        10'b 1001110111 :   address_offset = 12'b 100101110100 ;
        10'b 1001111000 :   address_offset = 12'b 100101111000 ;
        10'b 1001111001 :   address_offset = 12'b 100101111100 ;
        10'b 1001111010 :   address_offset = 12'b 100110000000 ;
        10'b 1001111011 :   address_offset = 12'b 100100010100 ;
        10'b 1001111100 :   address_offset = 12'b 100100011000 ;
        10'b 1001111101 :   address_offset = 12'b 100100011100 ;
        10'b 1001111110 :   address_offset = 12'b 100100100000 ;
        10'b 1001111111 :   address_offset = 12'b 100010110100 ;
        10'b 1010000000 :   address_offset = 12'b 100010111000 ;
        10'b 1010000001 :   address_offset = 12'b 100010111100 ;
        10'b 1010000010 :   address_offset = 12'b 000000000000 ;
        10'b 1010000011 :   address_offset = 12'b 000000000000 ;
        10'b 1010000100 :   address_offset = 12'b 101101101100 ;
        10'b 1010000101 :   address_offset = 12'b 101101110000 ;
        10'b 1010000110 :   address_offset = 12'b 101101110100 ;
        10'b 1010000111 :   address_offset = 12'b 101101111000 ;
        10'b 1010001000 :   address_offset = 12'b 101100001100 ;
        10'b 1010001001 :   address_offset = 12'b 101100010000 ;
        10'b 1010001010 :   address_offset = 12'b 101100010100 ;
        10'b 1010001011 :   address_offset = 12'b 101100011000 ;
        10'b 1010001100 :   address_offset = 12'b 101010101100 ;
        10'b 1010001101 :   address_offset = 12'b 101010101100 ;
        10'b 1010001110 :   address_offset = 12'b 101010110000 ;
        10'b 1010001111 :   address_offset = 12'b 101001000100 ;
        10'b 1010010000 :   address_offset = 12'b 101001001000 ;
        10'b 1010010001 :   address_offset = 12'b 101001001100 ;
        10'b 1010010010 :   address_offset = 12'b 101001010000 ;
        10'b 1010010011 :   address_offset = 12'b 100111100100 ;
        10'b 1010010100 :   address_offset = 12'b 100111101000 ;
        10'b 1010010101 :   address_offset = 12'b 100111101100 ;
        10'b 1010010110 :   address_offset = 12'b 100111110000 ;
        10'b 1010010111 :   address_offset = 12'b 100110000100 ;
        10'b 1010011000 :   address_offset = 12'b 100110001000 ;
        10'b 1010011001 :   address_offset = 12'b 100110001100 ;
        10'b 1010011010 :   address_offset = 12'b 100110010000 ;
        10'b 1010011011 :   address_offset = 12'b 100100100100 ;
        10'b 1010011100 :   address_offset = 12'b 100100101000 ;
        10'b 1010011101 :   address_offset = 12'b 100100101100 ;
        10'b 1010011110 :   address_offset = 12'b 000000000000 ;
        10'b 1010011111 :   address_offset = 12'b 000000000000 ;
        10'b 1010100000 :   address_offset = 12'b 101111011100 ;
        10'b 1010100001 :   address_offset = 12'b 101111100000 ;
        10'b 1010100010 :   address_offset = 12'b 101111100100 ;
        10'b 1010100011 :   address_offset = 12'b 101111101000 ;
        10'b 1010100100 :   address_offset = 12'b 101101111100 ;
        10'b 1010100101 :   address_offset = 12'b 101110000000 ;
        10'b 1010100110 :   address_offset = 12'b 101110000100 ;
        10'b 1010100111 :   address_offset = 12'b 101100011000 ;
        10'b 1010101000 :   address_offset = 12'b 101100011100 ;
        10'b 1010101001 :   address_offset = 12'b 101100100000 ;
        10'b 1010101010 :   address_offset = 12'b 101100100100 ;
        10'b 1010101011 :   address_offset = 12'b 101010111000 ;
        10'b 1010101100 :   address_offset = 12'b 101010111100 ;
        10'b 1010101101 :   address_offset = 12'b 101011000000 ;
        10'b 1010101110 :   address_offset = 12'b 101011000100 ;
        10'b 1010101111 :   address_offset = 12'b 101001011000 ;
        10'b 1010110000 :   address_offset = 12'b 101001011100 ;
        10'b 1010110001 :   address_offset = 12'b 101001011100 ;
        10'b 1010110010 :   address_offset = 12'b 101001100000 ;
        10'b 1010110011 :   address_offset = 12'b 100111110100 ;
        10'b 1010110100 :   address_offset = 12'b 100111111000 ;
        10'b 1010110101 :   address_offset = 12'b 100111111100 ;
        10'b 1010110110 :   address_offset = 12'b 101000000000 ;
        10'b 1010110111 :   address_offset = 12'b 100110010100 ;
        10'b 1010111000 :   address_offset = 12'b 100110011000 ;
        10'b 1010111001 :   address_offset = 12'b 100110011100 ;
        10'b 1010111010 :   address_offset = 12'b 000000000000 ;
        10'b 1010111011 :   address_offset = 12'b 000000000000 ;
        10'b 1010111100 :   address_offset = 12'b 000000000000 ;
        10'b 1010111101 :   address_offset = 12'b 000000000000 ;
        10'b 1010111110 :   address_offset = 12'b 000000000000 ;
        10'b 1010111111 :   address_offset = 12'b 101111101000 ;
        10'b 1011000000 :   address_offset = 12'b 101111101100 ;
        10'b 1011000001 :   address_offset = 12'b 101111110000 ;
        10'b 1011000010 :   address_offset = 12'b 101111110100 ;
        10'b 1011000011 :   address_offset = 12'b 101110001000 ;
        10'b 1011000100 :   address_offset = 12'b 101110001100 ;
        10'b 1011000101 :   address_offset = 12'b 101110010000 ;
        10'b 1011000110 :   address_offset = 12'b 101110010100 ;
        10'b 1011000111 :   address_offset = 12'b 101100101000 ;
        10'b 1011001000 :   address_offset = 12'b 101100101100 ;
        10'b 1011001001 :   address_offset = 12'b 101100110000 ;
        10'b 1011001010 :   address_offset = 12'b 101100110100 ;
        10'b 1011001011 :   address_offset = 12'b 101011001000 ;
        10'b 1011001100 :   address_offset = 12'b 101011001100 ;
        10'b 1011001101 :   address_offset = 12'b 101011010000 ;
        10'b 1011001110 :   address_offset = 12'b 101011010100 ;
        10'b 1011001111 :   address_offset = 12'b 101001101000 ;
        10'b 1011010000 :   address_offset = 12'b 101001101100 ;
        10'b 1011010001 :   address_offset = 12'b 101001110000 ;
        10'b 1011010010 :   address_offset = 12'b 101001110100 ;
        10'b 1011010011 :   address_offset = 12'b 101000001000 ;
        10'b 1011010100 :   address_offset = 12'b 101000001100 ;
        10'b 1011010101 :   address_offset = 12'b 101000001100 ;
        10'b 1011010110 :   address_offset = 12'b 000000000000 ;
        10'b 1011010111 :   address_offset = 12'b 000000000000 ;
        10'b 1011011000 :   address_offset = 12'b 000000000000 ;
        10'b 1011011001 :   address_offset = 12'b 000000000000 ;
        10'b 1011011010 :   address_offset = 12'b 000000000000 ;
        10'b 1011011011 :   address_offset = 12'b 000000000000 ;
        10'b 1011011100 :   address_offset = 12'b 000000000000 ;
        10'b 1011011101 :   address_offset = 12'b 000000000000 ;
        10'b 1011011110 :   address_offset = 12'b 000000000000 ;
        10'b 1011011111 :   address_offset = 12'b 101111111000 ;
        10'b 1011100000 :   address_offset = 12'b 101111111100 ;
        10'b 1011100001 :   address_offset = 12'b 110000000000 ;
        10'b 1011100010 :   address_offset = 12'b 110000000100 ;
        10'b 1011100011 :   address_offset = 12'b 101110011000 ;
        10'b 1011100100 :   address_offset = 12'b 101110011100 ;
        10'b 1011100101 :   address_offset = 12'b 101110100000 ;
        10'b 1011100110 :   address_offset = 12'b 101110100100 ;
        10'b 1011100111 :   address_offset = 12'b 101100111000 ;
        10'b 1011101000 :   address_offset = 12'b 101100111100 ;
        10'b 1011101001 :   address_offset = 12'b 101101000000 ;
        10'b 1011101010 :   address_offset = 12'b 101101000100 ;
        10'b 1011101011 :   address_offset = 12'b 101011011000 ;
        10'b 1011101100 :   address_offset = 12'b 101011011100 ;
        10'b 1011101101 :   address_offset = 12'b 101011100000 ;
        10'b 1011101110 :   address_offset = 12'b 101011100100 ;
        10'b 1011101111 :   address_offset = 12'b 101001111000 ;
        10'b 1011110000 :   address_offset = 12'b 101001111100 ;
        10'b 1011110001 :   address_offset = 12'b 000000000000 ;
        10'b 1011110010 :   address_offset = 12'b 000000000000 ;
        10'b 1011110011 :   address_offset = 12'b 000000000000 ;
        10'b 1011110100 :   address_offset = 12'b 000000000000 ;
        10'b 1011110101 :   address_offset = 12'b 000000000000 ;
        10'b 1011110110 :   address_offset = 12'b 000000000000 ;
        10'b 1011110111 :   address_offset = 12'b 000000000000 ;
        10'b 1011111000 :   address_offset = 12'b 000000000000 ;
        10'b 1011111001 :   address_offset = 12'b 000000000000 ;
        10'b 1011111010 :   address_offset = 12'b 000000000000 ;
        10'b 1011111011 :   address_offset = 12'b 000000000000 ;
        10'b 1011111100 :   address_offset = 12'b 000000000000 ;
        10'b 1011111101 :   address_offset = 12'b 000000000000 ;
        10'b 1011111110 :   address_offset = 12'b 000000000000 ;
        10'b 1011111111 :   address_offset = 12'b 110000001000 ;
        10'b 1100000000 :   address_offset = 12'b 110000001100 ;
        10'b 1100000001 :   address_offset = 12'b 110000010000 ;
        10'b 1100000010 :   address_offset = 12'b 110000010100 ;
        10'b 1100000011 :   address_offset = 12'b 101110101000 ;
        10'b 1100000100 :   address_offset = 12'b 101110101100 ;
        10'b 1100000101 :   address_offset = 12'b 101110110000 ;
        10'b 1100000110 :   address_offset = 12'b 101110110100 ;
        10'b 1100000111 :   address_offset = 12'b 101101001000 ;
        10'b 1100001000 :   address_offset = 12'b 101101001100 ;
        10'b 1100001001 :   address_offset = 12'b 101101010000 ;
        10'b 1100001010 :   address_offset = 12'b 101011100100 ;
        10'b 1100001011 :   address_offset = 12'b 101011101000 ;
        10'b 1100001100 :   address_offset = 12'b 101011101100 ;
        10'b 1100001101 :   address_offset = 12'b 000000000000 ;
        10'b 1100001110 :   address_offset = 12'b 000000000000 ;
        10'b 1100001111 :   address_offset = 12'b 000000000000 ;


        default: address_offset = 12'b0;
      endcase
    end 


endmodule
