module LUT_size16                                               // LUT to crop and resize, before resizing a dimension of 16 pixels
    (
        input logic [9:0] pixel_counter,                        // pixel number of the image after cropping
        output logic [9:0] address_offset                       // offset of the pixel value it should be stored in memory
    );
    
    logic [9:0] byte_offset;
    
    always_comb begin
        case (pixel_counter)
            10'b 0000000000 :   byte_offset = 10'b 0010101110;
            10'b 0000000001 :   byte_offset = 10'b 0010101111;
            10'b 0000000010 :   byte_offset = 10'b 0010101111;
            10'b 0000000011 :   byte_offset = 10'b 0010110000;
            10'b 0000000100 :   byte_offset = 10'b 0010110000;
            10'b 0000000101 :   byte_offset = 10'b 0010110001;
            10'b 0000000110 :   byte_offset = 10'b 0010110001;
            10'b 0000000111 :   byte_offset = 10'b 0010110010;
            10'b 0000001000 :   byte_offset = 10'b 0010110011;
            10'b 0000001001 :   byte_offset = 10'b 0010110011;
            10'b 0000001010 :   byte_offset = 10'b 0010110100;
            10'b 0000001011 :   byte_offset = 10'b 0010110100;
            10'b 0000001100 :   byte_offset = 10'b 0010110101;
            10'b 0000001101 :   byte_offset = 10'b 0010110101;
            10'b 0000001110 :   byte_offset = 10'b 0010110110;
            10'b 0000001111 :   byte_offset = 10'b 0010110111;
            10'b 0000010000 :   byte_offset = 10'b 0010110111;
            10'b 0000010001 :   byte_offset = 10'b 0010111000;
            10'b 0000010010 :   byte_offset = 10'b 0010111000;
            10'b 0000010011 :   byte_offset = 10'b 0010111001;
            10'b 0000010100 :   byte_offset = 10'b 0010111001;
            10'b 0000010101 :   byte_offset = 10'b 0010111010;
            10'b 0000010110 :   byte_offset = 10'b 0010111011;
            10'b 0000010111 :   byte_offset = 10'b 0010111011;
            10'b 0000011000 :   byte_offset = 10'b 0010111100;
            10'b 0000011001 :   byte_offset = 10'b 0010111100;
            10'b 0000011010 :   byte_offset = 10'b 0010111101;
            10'b 0000011011 :   byte_offset = 10'b 0010111101;
            10'b 0000011100 :   byte_offset = 10'b 0011001010;
            10'b 0000011101 :   byte_offset = 10'b 0011001011;
            10'b 0000011110 :   byte_offset = 10'b 0011001011;
            10'b 0000011111 :   byte_offset = 10'b 0011001100;
            10'b 0000100000 :   byte_offset = 10'b 0011001100;
            10'b 0000100001 :   byte_offset = 10'b 0011001101;
            10'b 0000100010 :   byte_offset = 10'b 0011001101;
            10'b 0000100011 :   byte_offset = 10'b 0011001110;
            10'b 0000100100 :   byte_offset = 10'b 0011001111;
            10'b 0000100101 :   byte_offset = 10'b 0011001111;
            10'b 0000100110 :   byte_offset = 10'b 0011010000;
            10'b 0000100111 :   byte_offset = 10'b 0011010000;
            10'b 0000101000 :   byte_offset = 10'b 0011010001;
            10'b 0000101001 :   byte_offset = 10'b 0011010001;
            10'b 0000101010 :   byte_offset = 10'b 0011010010;
            10'b 0000101011 :   byte_offset = 10'b 0011010011;
            10'b 0000101100 :   byte_offset = 10'b 0011010011;
            10'b 0000101101 :   byte_offset = 10'b 0011010100;
            10'b 0000101110 :   byte_offset = 10'b 0011010100;
            10'b 0000101111 :   byte_offset = 10'b 0011010101;
            10'b 0000110000 :   byte_offset = 10'b 0011010101;
            10'b 0000110001 :   byte_offset = 10'b 0011010110;
            10'b 0000110010 :   byte_offset = 10'b 0011010111;
            10'b 0000110011 :   byte_offset = 10'b 0011010111;
            10'b 0000110100 :   byte_offset = 10'b 0011011000;
            10'b 0000110101 :   byte_offset = 10'b 0011011000;
            10'b 0000110110 :   byte_offset = 10'b 0011011001;
            10'b 0000110111 :   byte_offset = 10'b 0011011001;
            10'b 0000111000 :   byte_offset = 10'b 0011001010;
            10'b 0000111001 :   byte_offset = 10'b 0011001011;
            10'b 0000111010 :   byte_offset = 10'b 0011001011;
            10'b 0000111011 :   byte_offset = 10'b 0011001100;
            10'b 0000111100 :   byte_offset = 10'b 0011001100;
            10'b 0000111101 :   byte_offset = 10'b 0011001101;
            10'b 0000111110 :   byte_offset = 10'b 0011001101;
            10'b 0000111111 :   byte_offset = 10'b 0011001110;
            10'b 0001000000 :   byte_offset = 10'b 0011001111;
            10'b 0001000001 :   byte_offset = 10'b 0011001111;
            10'b 0001000010 :   byte_offset = 10'b 0011010000;
            10'b 0001000011 :   byte_offset = 10'b 0011010000;
            10'b 0001000100 :   byte_offset = 10'b 0011010001;
            10'b 0001000101 :   byte_offset = 10'b 0011010001;
            10'b 0001000110 :   byte_offset = 10'b 0011010010;
            10'b 0001000111 :   byte_offset = 10'b 0011010011;
            10'b 0001001000 :   byte_offset = 10'b 0011010011;
            10'b 0001001001 :   byte_offset = 10'b 0011010100;
            10'b 0001001010 :   byte_offset = 10'b 0011010100;
            10'b 0001001011 :   byte_offset = 10'b 0011010101;
            10'b 0001001100 :   byte_offset = 10'b 0011010101;
            10'b 0001001101 :   byte_offset = 10'b 0011010110;
            10'b 0001001110 :   byte_offset = 10'b 0011010111;
            10'b 0001001111 :   byte_offset = 10'b 0011010111;
            10'b 0001010000 :   byte_offset = 10'b 0011011000;
            10'b 0001010001 :   byte_offset = 10'b 0011011000;
            10'b 0001010010 :   byte_offset = 10'b 0011011001;
            10'b 0001010011 :   byte_offset = 10'b 0011011001;
            10'b 0001010100 :   byte_offset = 10'b 0011100110;
            10'b 0001010101 :   byte_offset = 10'b 0011100111;
            10'b 0001010110 :   byte_offset = 10'b 0011100111;
            10'b 0001010111 :   byte_offset = 10'b 0011101000;
            10'b 0001011000 :   byte_offset = 10'b 0011101000;
            10'b 0001011001 :   byte_offset = 10'b 0011101001;
            10'b 0001011010 :   byte_offset = 10'b 0011101001;
            10'b 0001011011 :   byte_offset = 10'b 0011101010;
            10'b 0001011100 :   byte_offset = 10'b 0011101011;
            10'b 0001011101 :   byte_offset = 10'b 0011101011;
            10'b 0001011110 :   byte_offset = 10'b 0011101100;
            10'b 0001011111 :   byte_offset = 10'b 0011101100;
            10'b 0001100000 :   byte_offset = 10'b 0011101101;
            10'b 0001100001 :   byte_offset = 10'b 0011101101;
            10'b 0001100010 :   byte_offset = 10'b 0011101110;
            10'b 0001100011 :   byte_offset = 10'b 0011101111;
            10'b 0001100100 :   byte_offset = 10'b 0011101111;
            10'b 0001100101 :   byte_offset = 10'b 0011110000;
            10'b 0001100110 :   byte_offset = 10'b 0011110000;
            10'b 0001100111 :   byte_offset = 10'b 0011110001;
            10'b 0001101000 :   byte_offset = 10'b 0011110001;
            10'b 0001101001 :   byte_offset = 10'b 0011110010;
            10'b 0001101010 :   byte_offset = 10'b 0011110011;
            10'b 0001101011 :   byte_offset = 10'b 0011110011;
            10'b 0001101100 :   byte_offset = 10'b 0011110100;
            10'b 0001101101 :   byte_offset = 10'b 0011110100;
            10'b 0001101110 :   byte_offset = 10'b 0011110101;
            10'b 0001101111 :   byte_offset = 10'b 0011110101;
            10'b 0001110000 :   byte_offset = 10'b 0011100110;
            10'b 0001110001 :   byte_offset = 10'b 0011100111;
            10'b 0001110010 :   byte_offset = 10'b 0011100111;
            10'b 0001110011 :   byte_offset = 10'b 0011101000;
            10'b 0001110100 :   byte_offset = 10'b 0011101000;
            10'b 0001110101 :   byte_offset = 10'b 0011101001;
            10'b 0001110110 :   byte_offset = 10'b 0011101001;
            10'b 0001110111 :   byte_offset = 10'b 0011101010;
            10'b 0001111000 :   byte_offset = 10'b 0011101011;
            10'b 0001111001 :   byte_offset = 10'b 0011101011;
            10'b 0001111010 :   byte_offset = 10'b 0011101100;
            10'b 0001111011 :   byte_offset = 10'b 0011101100;
            10'b 0001111100 :   byte_offset = 10'b 0011101101;
            10'b 0001111101 :   byte_offset = 10'b 0011101101;
            10'b 0001111110 :   byte_offset = 10'b 0011101110;
            10'b 0001111111 :   byte_offset = 10'b 0011101111;
            10'b 0010000000 :   byte_offset = 10'b 0011101111;
            10'b 0010000001 :   byte_offset = 10'b 0011110000;
            10'b 0010000010 :   byte_offset = 10'b 0011110000;
            10'b 0010000011 :   byte_offset = 10'b 0011110001;
            10'b 0010000100 :   byte_offset = 10'b 0011110001;
            10'b 0010000101 :   byte_offset = 10'b 0011110010;
            10'b 0010000110 :   byte_offset = 10'b 0011110011;
            10'b 0010000111 :   byte_offset = 10'b 0011110011;
            10'b 0010001000 :   byte_offset = 10'b 0011110100;
            10'b 0010001001 :   byte_offset = 10'b 0011110100;
            10'b 0010001010 :   byte_offset = 10'b 0011110101;
            10'b 0010001011 :   byte_offset = 10'b 0011110101;
            10'b 0010001100 :   byte_offset = 10'b 0100000010;
            10'b 0010001101 :   byte_offset = 10'b 0100000011;
            10'b 0010001110 :   byte_offset = 10'b 0100000011;
            10'b 0010001111 :   byte_offset = 10'b 0100000100;
            10'b 0010010000 :   byte_offset = 10'b 0100000100;
            10'b 0010010001 :   byte_offset = 10'b 0100000101;
            10'b 0010010010 :   byte_offset = 10'b 0100000101;
            10'b 0010010011 :   byte_offset = 10'b 0100000110;
            10'b 0010010100 :   byte_offset = 10'b 0100000111;
            10'b 0010010101 :   byte_offset = 10'b 0100000111;
            10'b 0010010110 :   byte_offset = 10'b 0100001000;
            10'b 0010010111 :   byte_offset = 10'b 0100001000;
            10'b 0010011000 :   byte_offset = 10'b 0100001001;
            10'b 0010011001 :   byte_offset = 10'b 0100001001;
            10'b 0010011010 :   byte_offset = 10'b 0100001010;
            10'b 0010011011 :   byte_offset = 10'b 0100001011;
            10'b 0010011100 :   byte_offset = 10'b 0100001011;
            10'b 0010011101 :   byte_offset = 10'b 0100001100;
            10'b 0010011110 :   byte_offset = 10'b 0100001100;
            10'b 0010011111 :   byte_offset = 10'b 0100001101;
            10'b 0010100000 :   byte_offset = 10'b 0100001101;
            10'b 0010100001 :   byte_offset = 10'b 0100001110;
            10'b 0010100010 :   byte_offset = 10'b 0100001111;
            10'b 0010100011 :   byte_offset = 10'b 0100001111;
            10'b 0010100100 :   byte_offset = 10'b 0100010000;
            10'b 0010100101 :   byte_offset = 10'b 0100010000;
            10'b 0010100110 :   byte_offset = 10'b 0100010001;
            10'b 0010100111 :   byte_offset = 10'b 0100010001;
            10'b 0010101000 :   byte_offset = 10'b 0100000010;
            10'b 0010101001 :   byte_offset = 10'b 0100000011;
            10'b 0010101010 :   byte_offset = 10'b 0100000011;
            10'b 0010101011 :   byte_offset = 10'b 0100000100;
            10'b 0010101100 :   byte_offset = 10'b 0100000100;
            10'b 0010101101 :   byte_offset = 10'b 0100000101;
            10'b 0010101110 :   byte_offset = 10'b 0100000101;
            10'b 0010101111 :   byte_offset = 10'b 0100000110;
            10'b 0010110000 :   byte_offset = 10'b 0100000111;
            10'b 0010110001 :   byte_offset = 10'b 0100000111;
            10'b 0010110010 :   byte_offset = 10'b 0100001000;
            10'b 0010110011 :   byte_offset = 10'b 0100001000;
            10'b 0010110100 :   byte_offset = 10'b 0100001001;
            10'b 0010110101 :   byte_offset = 10'b 0100001001;
            10'b 0010110110 :   byte_offset = 10'b 0100001010;
            10'b 0010110111 :   byte_offset = 10'b 0100001011;
            10'b 0010111000 :   byte_offset = 10'b 0100001011;
            10'b 0010111001 :   byte_offset = 10'b 0100001100;
            10'b 0010111010 :   byte_offset = 10'b 0100001100;
            10'b 0010111011 :   byte_offset = 10'b 0100001101;
            10'b 0010111100 :   byte_offset = 10'b 0100001101;
            10'b 0010111101 :   byte_offset = 10'b 0100001110;
            10'b 0010111110 :   byte_offset = 10'b 0100001111;
            10'b 0010111111 :   byte_offset = 10'b 0100001111;
            10'b 0011000000 :   byte_offset = 10'b 0100010000;
            10'b 0011000001 :   byte_offset = 10'b 0100010000;
            10'b 0011000010 :   byte_offset = 10'b 0100010001;
            10'b 0011000011 :   byte_offset = 10'b 0100010001;
            10'b 0011000100 :   byte_offset = 10'b 0100011110;
            10'b 0011000101 :   byte_offset = 10'b 0100011111;
            10'b 0011000110 :   byte_offset = 10'b 0100011111;
            10'b 0011000111 :   byte_offset = 10'b 0100100000;
            10'b 0011001000 :   byte_offset = 10'b 0100100000;
            10'b 0011001001 :   byte_offset = 10'b 0100100001;
            10'b 0011001010 :   byte_offset = 10'b 0100100001;
            10'b 0011001011 :   byte_offset = 10'b 0100100010;
            10'b 0011001100 :   byte_offset = 10'b 0100100011;
            10'b 0011001101 :   byte_offset = 10'b 0100100011;
            10'b 0011001110 :   byte_offset = 10'b 0100100100;
            10'b 0011001111 :   byte_offset = 10'b 0100100100;
            10'b 0011010000 :   byte_offset = 10'b 0100100101;
            10'b 0011010001 :   byte_offset = 10'b 0100100101;
            10'b 0011010010 :   byte_offset = 10'b 0100100110;
            10'b 0011010011 :   byte_offset = 10'b 0100100111;
            10'b 0011010100 :   byte_offset = 10'b 0100100111;
            10'b 0011010101 :   byte_offset = 10'b 0100101000;
            10'b 0011010110 :   byte_offset = 10'b 0100101000;
            10'b 0011010111 :   byte_offset = 10'b 0100101001;
            10'b 0011011000 :   byte_offset = 10'b 0100101001;
            10'b 0011011001 :   byte_offset = 10'b 0100101010;
            10'b 0011011010 :   byte_offset = 10'b 0100101011;
            10'b 0011011011 :   byte_offset = 10'b 0100101011;
            10'b 0011011100 :   byte_offset = 10'b 0100101100;
            10'b 0011011101 :   byte_offset = 10'b 0100101100;
            10'b 0011011110 :   byte_offset = 10'b 0100101101;
            10'b 0011011111 :   byte_offset = 10'b 0100101101;
            10'b 0011100000 :   byte_offset = 10'b 0100111010;
            10'b 0011100001 :   byte_offset = 10'b 0100111011;
            10'b 0011100010 :   byte_offset = 10'b 0100111011;
            10'b 0011100011 :   byte_offset = 10'b 0100111100;
            10'b 0011100100 :   byte_offset = 10'b 0100111100;
            10'b 0011100101 :   byte_offset = 10'b 0100111101;
            10'b 0011100110 :   byte_offset = 10'b 0100111101;
            10'b 0011100111 :   byte_offset = 10'b 0100111110;
            10'b 0011101000 :   byte_offset = 10'b 0100111111;
            10'b 0011101001 :   byte_offset = 10'b 0100111111;
            10'b 0011101010 :   byte_offset = 10'b 0101000000;
            10'b 0011101011 :   byte_offset = 10'b 0101000000;
            10'b 0011101100 :   byte_offset = 10'b 0101000001;
            10'b 0011101101 :   byte_offset = 10'b 0101000001;
            10'b 0011101110 :   byte_offset = 10'b 0101000010;
            10'b 0011101111 :   byte_offset = 10'b 0101000011;
            10'b 0011110000 :   byte_offset = 10'b 0101000011;
            10'b 0011110001 :   byte_offset = 10'b 0101000100;
            10'b 0011110010 :   byte_offset = 10'b 0101000100;
            10'b 0011110011 :   byte_offset = 10'b 0101000101;
            10'b 0011110100 :   byte_offset = 10'b 0101000101;
            10'b 0011110101 :   byte_offset = 10'b 0101000110;
            10'b 0011110110 :   byte_offset = 10'b 0101000111;
            10'b 0011110111 :   byte_offset = 10'b 0101000111;
            10'b 0011111000 :   byte_offset = 10'b 0101001000;
            10'b 0011111001 :   byte_offset = 10'b 0101001000;
            10'b 0011111010 :   byte_offset = 10'b 0101001001;
            10'b 0011111011 :   byte_offset = 10'b 0101001001;
            10'b 0011111100 :   byte_offset = 10'b 0100111010;
            10'b 0011111101 :   byte_offset = 10'b 0100111011;
            10'b 0011111110 :   byte_offset = 10'b 0100111011;
            10'b 0011111111 :   byte_offset = 10'b 0100111100;
            10'b 0100000000 :   byte_offset = 10'b 0100111100;
            10'b 0100000001 :   byte_offset = 10'b 0100111101;
            10'b 0100000010 :   byte_offset = 10'b 0100111101;
            10'b 0100000011 :   byte_offset = 10'b 0100111110;
            10'b 0100000100 :   byte_offset = 10'b 0100111111;
            10'b 0100000101 :   byte_offset = 10'b 0100111111;
            10'b 0100000110 :   byte_offset = 10'b 0101000000;
            10'b 0100000111 :   byte_offset = 10'b 0101000000;
            10'b 0100001000 :   byte_offset = 10'b 0101000001;
            10'b 0100001001 :   byte_offset = 10'b 0101000001;
            10'b 0100001010 :   byte_offset = 10'b 0101000010;
            10'b 0100001011 :   byte_offset = 10'b 0101000011;
            10'b 0100001100 :   byte_offset = 10'b 0101000011;
            10'b 0100001101 :   byte_offset = 10'b 0101000100;
            10'b 0100001110 :   byte_offset = 10'b 0101000100;
            10'b 0100001111 :   byte_offset = 10'b 0101000101;
            10'b 0100010000 :   byte_offset = 10'b 0101000101;
            10'b 0100010001 :   byte_offset = 10'b 0101000110;
            10'b 0100010010 :   byte_offset = 10'b 0101000111;
            10'b 0100010011 :   byte_offset = 10'b 0101000111;
            10'b 0100010100 :   byte_offset = 10'b 0101001000;
            10'b 0100010101 :   byte_offset = 10'b 0101001000;
            10'b 0100010110 :   byte_offset = 10'b 0101001001;
            10'b 0100010111 :   byte_offset = 10'b 0101001001;
            10'b 0100011000 :   byte_offset = 10'b 0101010110;
            10'b 0100011001 :   byte_offset = 10'b 0101010111;
            10'b 0100011010 :   byte_offset = 10'b 0101010111;
            10'b 0100011011 :   byte_offset = 10'b 0101011000;
            10'b 0100011100 :   byte_offset = 10'b 0101011000;
            10'b 0100011101 :   byte_offset = 10'b 0101011001;
            10'b 0100011110 :   byte_offset = 10'b 0101011001;
            10'b 0100011111 :   byte_offset = 10'b 0101011010;
            10'b 0100100000 :   byte_offset = 10'b 0101011011;
            10'b 0100100001 :   byte_offset = 10'b 0101011011;
            10'b 0100100010 :   byte_offset = 10'b 0101011100;
            10'b 0100100011 :   byte_offset = 10'b 0101011100;
            10'b 0100100100 :   byte_offset = 10'b 0101011101;
            10'b 0100100101 :   byte_offset = 10'b 0101011101;
            10'b 0100100110 :   byte_offset = 10'b 0101011110;
            10'b 0100100111 :   byte_offset = 10'b 0101011111;
            10'b 0100101000 :   byte_offset = 10'b 0101011111;
            10'b 0100101001 :   byte_offset = 10'b 0101100000;
            10'b 0100101010 :   byte_offset = 10'b 0101100000;
            10'b 0100101011 :   byte_offset = 10'b 0101100001;
            10'b 0100101100 :   byte_offset = 10'b 0101100001;
            10'b 0100101101 :   byte_offset = 10'b 0101100010;
            10'b 0100101110 :   byte_offset = 10'b 0101100011;
            10'b 0100101111 :   byte_offset = 10'b 0101100011;
            10'b 0100110000 :   byte_offset = 10'b 0101100100;
            10'b 0100110001 :   byte_offset = 10'b 0101100100;
            10'b 0100110010 :   byte_offset = 10'b 0101100101;
            10'b 0100110011 :   byte_offset = 10'b 0101100101;
            10'b 0100110100 :   byte_offset = 10'b 0101010110;
            10'b 0100110101 :   byte_offset = 10'b 0101010111;
            10'b 0100110110 :   byte_offset = 10'b 0101010111;
            10'b 0100110111 :   byte_offset = 10'b 0101011000;
            10'b 0100111000 :   byte_offset = 10'b 0101011000;
            10'b 0100111001 :   byte_offset = 10'b 0101011001;
            10'b 0100111010 :   byte_offset = 10'b 0101011001;
            10'b 0100111011 :   byte_offset = 10'b 0101011010;
            10'b 0100111100 :   byte_offset = 10'b 0101011011;
            10'b 0100111101 :   byte_offset = 10'b 0101011011;
            10'b 0100111110 :   byte_offset = 10'b 0101011100;
            10'b 0100111111 :   byte_offset = 10'b 0101011100;
            10'b 0101000000 :   byte_offset = 10'b 0101011101;
            10'b 0101000001 :   byte_offset = 10'b 0101011101;
            10'b 0101000010 :   byte_offset = 10'b 0101011110;
            10'b 0101000011 :   byte_offset = 10'b 0101011111;
            10'b 0101000100 :   byte_offset = 10'b 0101011111;
            10'b 0101000101 :   byte_offset = 10'b 0101100000;
            10'b 0101000110 :   byte_offset = 10'b 0101100000;
            10'b 0101000111 :   byte_offset = 10'b 0101100001;
            10'b 0101001000 :   byte_offset = 10'b 0101100001;
            10'b 0101001001 :   byte_offset = 10'b 0101100010;
            10'b 0101001010 :   byte_offset = 10'b 0101100011;
            10'b 0101001011 :   byte_offset = 10'b 0101100011;
            10'b 0101001100 :   byte_offset = 10'b 0101100100;
            10'b 0101001101 :   byte_offset = 10'b 0101100100;
            10'b 0101001110 :   byte_offset = 10'b 0101100101;
            10'b 0101001111 :   byte_offset = 10'b 0101100101;
            10'b 0101010000 :   byte_offset = 10'b 0101110010;
            10'b 0101010001 :   byte_offset = 10'b 0101110011;
            10'b 0101010010 :   byte_offset = 10'b 0101110011;
            10'b 0101010011 :   byte_offset = 10'b 0101110100;
            10'b 0101010100 :   byte_offset = 10'b 0101110100;
            10'b 0101010101 :   byte_offset = 10'b 0101110101;
            10'b 0101010110 :   byte_offset = 10'b 0101110101;
            10'b 0101010111 :   byte_offset = 10'b 0101110110;
            10'b 0101011000 :   byte_offset = 10'b 0101110111;
            10'b 0101011001 :   byte_offset = 10'b 0101110111;
            10'b 0101011010 :   byte_offset = 10'b 0101111000;
            10'b 0101011011 :   byte_offset = 10'b 0101111000;
            10'b 0101011100 :   byte_offset = 10'b 0101111001;
            10'b 0101011101 :   byte_offset = 10'b 0101111001;
            10'b 0101011110 :   byte_offset = 10'b 0101111010;
            10'b 0101011111 :   byte_offset = 10'b 0101111011;
            10'b 0101100000 :   byte_offset = 10'b 0101111011;
            10'b 0101100001 :   byte_offset = 10'b 0101111100;
            10'b 0101100010 :   byte_offset = 10'b 0101111100;
            10'b 0101100011 :   byte_offset = 10'b 0101111101;
            10'b 0101100100 :   byte_offset = 10'b 0101111101;
            10'b 0101100101 :   byte_offset = 10'b 0101111110;
            10'b 0101100110 :   byte_offset = 10'b 0101111111;
            10'b 0101100111 :   byte_offset = 10'b 0101111111;
            10'b 0101101000 :   byte_offset = 10'b 0110000000;
            10'b 0101101001 :   byte_offset = 10'b 0110000000;
            10'b 0101101010 :   byte_offset = 10'b 0110000001;
            10'b 0101101011 :   byte_offset = 10'b 0110000001;
            10'b 0101101100 :   byte_offset = 10'b 0101110010;
            10'b 0101101101 :   byte_offset = 10'b 0101110011;
            10'b 0101101110 :   byte_offset = 10'b 0101110011;
            10'b 0101101111 :   byte_offset = 10'b 0101110100;
            10'b 0101110000 :   byte_offset = 10'b 0101110100;
            10'b 0101110001 :   byte_offset = 10'b 0101110101;
            10'b 0101110010 :   byte_offset = 10'b 0101110101;
            10'b 0101110011 :   byte_offset = 10'b 0101110110;
            10'b 0101110100 :   byte_offset = 10'b 0101110111;
            10'b 0101110101 :   byte_offset = 10'b 0101110111;
            10'b 0101110110 :   byte_offset = 10'b 0101111000;
            10'b 0101110111 :   byte_offset = 10'b 0101111000;
            10'b 0101111000 :   byte_offset = 10'b 0101111001;
            10'b 0101111001 :   byte_offset = 10'b 0101111001;
            10'b 0101111010 :   byte_offset = 10'b 0101111010;
            10'b 0101111011 :   byte_offset = 10'b 0101111011;
            10'b 0101111100 :   byte_offset = 10'b 0101111011;
            10'b 0101111101 :   byte_offset = 10'b 0101111100;
            10'b 0101111110 :   byte_offset = 10'b 0101111100;
            10'b 0101111111 :   byte_offset = 10'b 0101111101;
            10'b 0110000000 :   byte_offset = 10'b 0101111101;
            10'b 0110000001 :   byte_offset = 10'b 0101111110;
            10'b 0110000010 :   byte_offset = 10'b 0101111111;
            10'b 0110000011 :   byte_offset = 10'b 0101111111;
            10'b 0110000100 :   byte_offset = 10'b 0110000000;
            10'b 0110000101 :   byte_offset = 10'b 0110000000;
            10'b 0110000110 :   byte_offset = 10'b 0110000001;
            10'b 0110000111 :   byte_offset = 10'b 0110000001;
            10'b 0110001000 :   byte_offset = 10'b 0110001110;
            10'b 0110001001 :   byte_offset = 10'b 0110001111;
            10'b 0110001010 :   byte_offset = 10'b 0110001111;
            10'b 0110001011 :   byte_offset = 10'b 0110010000;
            10'b 0110001100 :   byte_offset = 10'b 0110010000;
            10'b 0110001101 :   byte_offset = 10'b 0110010001;
            10'b 0110001110 :   byte_offset = 10'b 0110010001;
            10'b 0110001111 :   byte_offset = 10'b 0110010010;
            10'b 0110010000 :   byte_offset = 10'b 0110010011;
            10'b 0110010001 :   byte_offset = 10'b 0110010011;
            10'b 0110010010 :   byte_offset = 10'b 0110010100;
            10'b 0110010011 :   byte_offset = 10'b 0110010100;
            10'b 0110010100 :   byte_offset = 10'b 0110010101;
            10'b 0110010101 :   byte_offset = 10'b 0110010101;
            10'b 0110010110 :   byte_offset = 10'b 0110010110;
            10'b 0110010111 :   byte_offset = 10'b 0110010111;
            10'b 0110011000 :   byte_offset = 10'b 0110010111;
            10'b 0110011001 :   byte_offset = 10'b 0110011000;
            10'b 0110011010 :   byte_offset = 10'b 0110011000;
            10'b 0110011011 :   byte_offset = 10'b 0110011001;
            10'b 0110011100 :   byte_offset = 10'b 0110011001;
            10'b 0110011101 :   byte_offset = 10'b 0110011010;
            10'b 0110011110 :   byte_offset = 10'b 0110011011;
            10'b 0110011111 :   byte_offset = 10'b 0110011011;
            10'b 0110100000 :   byte_offset = 10'b 0110011100;
            10'b 0110100001 :   byte_offset = 10'b 0110011100;
            10'b 0110100010 :   byte_offset = 10'b 0110011101;
            10'b 0110100011 :   byte_offset = 10'b 0110011101;
            10'b 0110100100 :   byte_offset = 10'b 0110101010;
            10'b 0110100101 :   byte_offset = 10'b 0110101011;
            10'b 0110100110 :   byte_offset = 10'b 0110101011;
            10'b 0110100111 :   byte_offset = 10'b 0110101100;
            10'b 0110101000 :   byte_offset = 10'b 0110101100;
            10'b 0110101001 :   byte_offset = 10'b 0110101101;
            10'b 0110101010 :   byte_offset = 10'b 0110101101;
            10'b 0110101011 :   byte_offset = 10'b 0110101110;
            10'b 0110101100 :   byte_offset = 10'b 0110101111;
            10'b 0110101101 :   byte_offset = 10'b 0110101111;
            10'b 0110101110 :   byte_offset = 10'b 0110110000;
            10'b 0110101111 :   byte_offset = 10'b 0110110000;
            10'b 0110110000 :   byte_offset = 10'b 0110110001;
            10'b 0110110001 :   byte_offset = 10'b 0110110001;
            10'b 0110110010 :   byte_offset = 10'b 0110110010;
            10'b 0110110011 :   byte_offset = 10'b 0110110011;
            10'b 0110110100 :   byte_offset = 10'b 0110110011;
            10'b 0110110101 :   byte_offset = 10'b 0110110100;
            10'b 0110110110 :   byte_offset = 10'b 0110110100;
            10'b 0110110111 :   byte_offset = 10'b 0110110101;
            10'b 0110111000 :   byte_offset = 10'b 0110110101;
            10'b 0110111001 :   byte_offset = 10'b 0110110110;
            10'b 0110111010 :   byte_offset = 10'b 0110110111;
            10'b 0110111011 :   byte_offset = 10'b 0110110111;
            10'b 0110111100 :   byte_offset = 10'b 0110111000;
            10'b 0110111101 :   byte_offset = 10'b 0110111000;
            10'b 0110111110 :   byte_offset = 10'b 0110111001;
            10'b 0110111111 :   byte_offset = 10'b 0110111001;
            10'b 0111000000 :   byte_offset = 10'b 0110101010;
            10'b 0111000001 :   byte_offset = 10'b 0110101011;
            10'b 0111000010 :   byte_offset = 10'b 0110101011;
            10'b 0111000011 :   byte_offset = 10'b 0110101100;
            10'b 0111000100 :   byte_offset = 10'b 0110101100;
            10'b 0111000101 :   byte_offset = 10'b 0110101101;
            10'b 0111000110 :   byte_offset = 10'b 0110101101;
            10'b 0111000111 :   byte_offset = 10'b 0110101110;
            10'b 0111001000 :   byte_offset = 10'b 0110101111;
            10'b 0111001001 :   byte_offset = 10'b 0110101111;
            10'b 0111001010 :   byte_offset = 10'b 0110110000;
            10'b 0111001011 :   byte_offset = 10'b 0110110000;
            10'b 0111001100 :   byte_offset = 10'b 0110110001;
            10'b 0111001101 :   byte_offset = 10'b 0110110001;
            10'b 0111001110 :   byte_offset = 10'b 0110110010;
            10'b 0111001111 :   byte_offset = 10'b 0110110011;
            10'b 0111010000 :   byte_offset = 10'b 0110110011;
            10'b 0111010001 :   byte_offset = 10'b 0110110100;
            10'b 0111010010 :   byte_offset = 10'b 0110110100;
            10'b 0111010011 :   byte_offset = 10'b 0110110101;
            10'b 0111010100 :   byte_offset = 10'b 0110110101;
            10'b 0111010101 :   byte_offset = 10'b 0110110110;
            10'b 0111010110 :   byte_offset = 10'b 0110110111;
            10'b 0111010111 :   byte_offset = 10'b 0110110111;
            10'b 0111011000 :   byte_offset = 10'b 0110111000;
            10'b 0111011001 :   byte_offset = 10'b 0110111000;
            10'b 0111011010 :   byte_offset = 10'b 0110111001;
            10'b 0111011011 :   byte_offset = 10'b 0110111001;
            10'b 0111011100 :   byte_offset = 10'b 0111000110;
            10'b 0111011101 :   byte_offset = 10'b 0111000111;
            10'b 0111011110 :   byte_offset = 10'b 0111000111;
            10'b 0111011111 :   byte_offset = 10'b 0111001000;
            10'b 0111100000 :   byte_offset = 10'b 0111001000;
            10'b 0111100001 :   byte_offset = 10'b 0111001001;
            10'b 0111100010 :   byte_offset = 10'b 0111001001;
            10'b 0111100011 :   byte_offset = 10'b 0111001010;
            10'b 0111100100 :   byte_offset = 10'b 0111001011;
            10'b 0111100101 :   byte_offset = 10'b 0111001011;
            10'b 0111100110 :   byte_offset = 10'b 0111001100;
            10'b 0111100111 :   byte_offset = 10'b 0111001100;
            10'b 0111101000 :   byte_offset = 10'b 0111001101;
            10'b 0111101001 :   byte_offset = 10'b 0111001101;
            10'b 0111101010 :   byte_offset = 10'b 0111001110;
            10'b 0111101011 :   byte_offset = 10'b 0111001111;
            10'b 0111101100 :   byte_offset = 10'b 0111001111;
            10'b 0111101101 :   byte_offset = 10'b 0111010000;
            10'b 0111101110 :   byte_offset = 10'b 0111010000;
            10'b 0111101111 :   byte_offset = 10'b 0111010001;
            10'b 0111110000 :   byte_offset = 10'b 0111010001;
            10'b 0111110001 :   byte_offset = 10'b 0111010010;
            10'b 0111110010 :   byte_offset = 10'b 0111010011;
            10'b 0111110011 :   byte_offset = 10'b 0111010011;
            10'b 0111110100 :   byte_offset = 10'b 0111010100;
            10'b 0111110101 :   byte_offset = 10'b 0111010100;
            10'b 0111110110 :   byte_offset = 10'b 0111010101;
            10'b 0111110111 :   byte_offset = 10'b 0111010101;
            10'b 0111111000 :   byte_offset = 10'b 0111000110;
            10'b 0111111001 :   byte_offset = 10'b 0111000111;
            10'b 0111111010 :   byte_offset = 10'b 0111000111;
            10'b 0111111011 :   byte_offset = 10'b 0111001000;
            10'b 0111111100 :   byte_offset = 10'b 0111001000;
            10'b 0111111101 :   byte_offset = 10'b 0111001001;
            10'b 0111111110 :   byte_offset = 10'b 0111001001;
            10'b 0111111111 :   byte_offset = 10'b 0111001010;
            10'b 1000000000 :   byte_offset = 10'b 0111001011;
            10'b 1000000001 :   byte_offset = 10'b 0111001011;
            10'b 1000000010 :   byte_offset = 10'b 0111001100;
            10'b 1000000011 :   byte_offset = 10'b 0111001100;
            10'b 1000000100 :   byte_offset = 10'b 0111001101;
            10'b 1000000101 :   byte_offset = 10'b 0111001101;
            10'b 1000000110 :   byte_offset = 10'b 0111001110;
            10'b 1000000111 :   byte_offset = 10'b 0111001111;
            10'b 1000001000 :   byte_offset = 10'b 0111001111;
            10'b 1000001001 :   byte_offset = 10'b 0111010000;
            10'b 1000001010 :   byte_offset = 10'b 0111010000;
            10'b 1000001011 :   byte_offset = 10'b 0111010001;
            10'b 1000001100 :   byte_offset = 10'b 0111010001;
            10'b 1000001101 :   byte_offset = 10'b 0111010010;
            10'b 1000001110 :   byte_offset = 10'b 0111010011;
            10'b 1000001111 :   byte_offset = 10'b 0111010011;
            10'b 1000010000 :   byte_offset = 10'b 0111010100;
            10'b 1000010001 :   byte_offset = 10'b 0111010100;
            10'b 1000010010 :   byte_offset = 10'b 0111010101;
            10'b 1000010011 :   byte_offset = 10'b 0111010101;
            10'b 1000010100 :   byte_offset = 10'b 0111100010;
            10'b 1000010101 :   byte_offset = 10'b 0111100011;
            10'b 1000010110 :   byte_offset = 10'b 0111100011;
            10'b 1000010111 :   byte_offset = 10'b 0111100100;
            10'b 1000011000 :   byte_offset = 10'b 0111100100;
            10'b 1000011001 :   byte_offset = 10'b 0111100101;
            10'b 1000011010 :   byte_offset = 10'b 0111100101;
            10'b 1000011011 :   byte_offset = 10'b 0111100110;
            10'b 1000011100 :   byte_offset = 10'b 0111100111;
            10'b 1000011101 :   byte_offset = 10'b 0111100111;
            10'b 1000011110 :   byte_offset = 10'b 0111101000;
            10'b 1000011111 :   byte_offset = 10'b 0111101000;
            10'b 1000100000 :   byte_offset = 10'b 0111101001;
            10'b 1000100001 :   byte_offset = 10'b 0111101001;
            10'b 1000100010 :   byte_offset = 10'b 0111101010;
            10'b 1000100011 :   byte_offset = 10'b 0111101011;
            10'b 1000100100 :   byte_offset = 10'b 0111101011;
            10'b 1000100101 :   byte_offset = 10'b 0111101100;
            10'b 1000100110 :   byte_offset = 10'b 0111101100;
            10'b 1000100111 :   byte_offset = 10'b 0111101101;
            10'b 1000101000 :   byte_offset = 10'b 0111101101;
            10'b 1000101001 :   byte_offset = 10'b 0111101110;
            10'b 1000101010 :   byte_offset = 10'b 0111101111;
            10'b 1000101011 :   byte_offset = 10'b 0111101111;
            10'b 1000101100 :   byte_offset = 10'b 0111110000;
            10'b 1000101101 :   byte_offset = 10'b 0111110000;
            10'b 1000101110 :   byte_offset = 10'b 0111110001;
            10'b 1000101111 :   byte_offset = 10'b 0111110001;
            10'b 1000110000 :   byte_offset = 10'b 0111100010;
            10'b 1000110001 :   byte_offset = 10'b 0111100011;
            10'b 1000110010 :   byte_offset = 10'b 0111100011;
            10'b 1000110011 :   byte_offset = 10'b 0111100100;
            10'b 1000110100 :   byte_offset = 10'b 0111100100;
            10'b 1000110101 :   byte_offset = 10'b 0111100101;
            10'b 1000110110 :   byte_offset = 10'b 0111100101;
            10'b 1000110111 :   byte_offset = 10'b 0111100110;
            10'b 1000111000 :   byte_offset = 10'b 0111100111;
            10'b 1000111001 :   byte_offset = 10'b 0111100111;
            10'b 1000111010 :   byte_offset = 10'b 0111101000;
            10'b 1000111011 :   byte_offset = 10'b 0111101000;
            10'b 1000111100 :   byte_offset = 10'b 0111101001;
            10'b 1000111101 :   byte_offset = 10'b 0111101001;
            10'b 1000111110 :   byte_offset = 10'b 0111101010;
            10'b 1000111111 :   byte_offset = 10'b 0111101011;
            10'b 1001000000 :   byte_offset = 10'b 0111101011;
            10'b 1001000001 :   byte_offset = 10'b 0111101100;
            10'b 1001000010 :   byte_offset = 10'b 0111101100;
            10'b 1001000011 :   byte_offset = 10'b 0111101101;
            10'b 1001000100 :   byte_offset = 10'b 0111101101;
            10'b 1001000101 :   byte_offset = 10'b 0111101110;
            10'b 1001000110 :   byte_offset = 10'b 0111101111;
            10'b 1001000111 :   byte_offset = 10'b 0111101111;
            10'b 1001001000 :   byte_offset = 10'b 0111110000;
            10'b 1001001001 :   byte_offset = 10'b 0111110000;
            10'b 1001001010 :   byte_offset = 10'b 0111110001;
            10'b 1001001011 :   byte_offset = 10'b 0111110001;
            10'b 1001001100 :   byte_offset = 10'b 0111111110;
            10'b 1001001101 :   byte_offset = 10'b 0111111111;
            10'b 1001001110 :   byte_offset = 10'b 0111111111;
            10'b 1001001111 :   byte_offset = 10'b 1000000000;
            10'b 1001010000 :   byte_offset = 10'b 1000000000;
            10'b 1001010001 :   byte_offset = 10'b 1000000001;
            10'b 1001010010 :   byte_offset = 10'b 1000000001;
            10'b 1001010011 :   byte_offset = 10'b 1000000010;
            10'b 1001010100 :   byte_offset = 10'b 1000000011;
            10'b 1001010101 :   byte_offset = 10'b 1000000011;
            10'b 1001010110 :   byte_offset = 10'b 1000000100;
            10'b 1001010111 :   byte_offset = 10'b 1000000100;
            10'b 1001011000 :   byte_offset = 10'b 1000000101;
            10'b 1001011001 :   byte_offset = 10'b 1000000101;
            10'b 1001011010 :   byte_offset = 10'b 1000000110;
            10'b 1001011011 :   byte_offset = 10'b 1000000111;
            10'b 1001011100 :   byte_offset = 10'b 1000000111;
            10'b 1001011101 :   byte_offset = 10'b 1000001000;
            10'b 1001011110 :   byte_offset = 10'b 1000001000;
            10'b 1001011111 :   byte_offset = 10'b 1000001001;
            10'b 1001100000 :   byte_offset = 10'b 1000001001;
            10'b 1001100001 :   byte_offset = 10'b 1000001010;
            10'b 1001100010 :   byte_offset = 10'b 1000001011;
            10'b 1001100011 :   byte_offset = 10'b 1000001011;
            10'b 1001100100 :   byte_offset = 10'b 1000001100;
            10'b 1001100101 :   byte_offset = 10'b 1000001100;
            10'b 1001100110 :   byte_offset = 10'b 1000001101;
            10'b 1001100111 :   byte_offset = 10'b 1000001101;
            10'b 1001101000 :   byte_offset = 10'b 1000011010;
            10'b 1001101001 :   byte_offset = 10'b 1000011011;
            10'b 1001101010 :   byte_offset = 10'b 1000011011;
            10'b 1001101011 :   byte_offset = 10'b 1000011100;
            10'b 1001101100 :   byte_offset = 10'b 1000011100;
            10'b 1001101101 :   byte_offset = 10'b 1000011101;
            10'b 1001101110 :   byte_offset = 10'b 1000011101;
            10'b 1001101111 :   byte_offset = 10'b 1000011110;
            10'b 1001110000 :   byte_offset = 10'b 1000011111;
            10'b 1001110001 :   byte_offset = 10'b 1000011111;
            10'b 1001110010 :   byte_offset = 10'b 1000100000;
            10'b 1001110011 :   byte_offset = 10'b 1000100000;
            10'b 1001110100 :   byte_offset = 10'b 1000100001;
            10'b 1001110101 :   byte_offset = 10'b 1000100001;
            10'b 1001110110 :   byte_offset = 10'b 1000100010;
            10'b 1001110111 :   byte_offset = 10'b 1000100011;
            10'b 1001111000 :   byte_offset = 10'b 1000100011;
            10'b 1001111001 :   byte_offset = 10'b 1000100100;
            10'b 1001111010 :   byte_offset = 10'b 1000100100;
            10'b 1001111011 :   byte_offset = 10'b 1000100101;
            10'b 1001111100 :   byte_offset = 10'b 1000100101;
            10'b 1001111101 :   byte_offset = 10'b 1000100110;
            10'b 1001111110 :   byte_offset = 10'b 1000100111;
            10'b 1001111111 :   byte_offset = 10'b 1000100111;
            10'b 1010000000 :   byte_offset = 10'b 1000101000;
            10'b 1010000001 :   byte_offset = 10'b 1000101000;
            10'b 1010000010 :   byte_offset = 10'b 1000101001;
            10'b 1010000011 :   byte_offset = 10'b 1000101001;
            10'b 1010000100 :   byte_offset = 10'b 1000011010;
            10'b 1010000101 :   byte_offset = 10'b 1000011011;
            10'b 1010000110 :   byte_offset = 10'b 1000011011;
            10'b 1010000111 :   byte_offset = 10'b 1000011100;
            10'b 1010001000 :   byte_offset = 10'b 1000011100;
            10'b 1010001001 :   byte_offset = 10'b 1000011101;
            10'b 1010001010 :   byte_offset = 10'b 1000011101;
            10'b 1010001011 :   byte_offset = 10'b 1000011110;
            10'b 1010001100 :   byte_offset = 10'b 1000011111;
            10'b 1010001101 :   byte_offset = 10'b 1000011111;
            10'b 1010001110 :   byte_offset = 10'b 1000100000;
            10'b 1010001111 :   byte_offset = 10'b 1000100000;
            10'b 1010010000 :   byte_offset = 10'b 1000100001;
            10'b 1010010001 :   byte_offset = 10'b 1000100001;
            10'b 1010010010 :   byte_offset = 10'b 1000100010;
            10'b 1010010011 :   byte_offset = 10'b 1000100011;
            10'b 1010010100 :   byte_offset = 10'b 1000100011;
            10'b 1010010101 :   byte_offset = 10'b 1000100100;
            10'b 1010010110 :   byte_offset = 10'b 1000100100;
            10'b 1010010111 :   byte_offset = 10'b 1000100101;
            10'b 1010011000 :   byte_offset = 10'b 1000100101;
            10'b 1010011001 :   byte_offset = 10'b 1000100110;
            10'b 1010011010 :   byte_offset = 10'b 1000100111;
            10'b 1010011011 :   byte_offset = 10'b 1000100111;
            10'b 1010011100 :   byte_offset = 10'b 1000101000;
            10'b 1010011101 :   byte_offset = 10'b 1000101000;
            10'b 1010011110 :   byte_offset = 10'b 1000101001;
            10'b 1010011111 :   byte_offset = 10'b 1000101001;
            10'b 1010100000 :   byte_offset = 10'b 1000110110;
            10'b 1010100001 :   byte_offset = 10'b 1000110111;
            10'b 1010100010 :   byte_offset = 10'b 1000110111;
            10'b 1010100011 :   byte_offset = 10'b 1000111000;
            10'b 1010100100 :   byte_offset = 10'b 1000111000;
            10'b 1010100101 :   byte_offset = 10'b 1000111001;
            10'b 1010100110 :   byte_offset = 10'b 1000111001;
            10'b 1010100111 :   byte_offset = 10'b 1000111010;
            10'b 1010101000 :   byte_offset = 10'b 1000111011;
            10'b 1010101001 :   byte_offset = 10'b 1000111011;
            10'b 1010101010 :   byte_offset = 10'b 1000111100;
            10'b 1010101011 :   byte_offset = 10'b 1000111100;
            10'b 1010101100 :   byte_offset = 10'b 1000111101;
            10'b 1010101101 :   byte_offset = 10'b 1000111101;
            10'b 1010101110 :   byte_offset = 10'b 1000111110;
            10'b 1010101111 :   byte_offset = 10'b 1000111111;
            10'b 1010110000 :   byte_offset = 10'b 1000111111;
            10'b 1010110001 :   byte_offset = 10'b 1001000000;
            10'b 1010110010 :   byte_offset = 10'b 1001000000;
            10'b 1010110011 :   byte_offset = 10'b 1001000001;
            10'b 1010110100 :   byte_offset = 10'b 1001000001;
            10'b 1010110101 :   byte_offset = 10'b 1001000010;
            10'b 1010110110 :   byte_offset = 10'b 1001000011;
            10'b 1010110111 :   byte_offset = 10'b 1001000011;
            10'b 1010111000 :   byte_offset = 10'b 1001000100;
            10'b 1010111001 :   byte_offset = 10'b 1001000100;
            10'b 1010111010 :   byte_offset = 10'b 1001000101;
            10'b 1010111011 :   byte_offset = 10'b 1001000101;
            10'b 1010111100 :   byte_offset = 10'b 1000110110;
            10'b 1010111101 :   byte_offset = 10'b 1000110111;
            10'b 1010111110 :   byte_offset = 10'b 1000110111;
            10'b 1010111111 :   byte_offset = 10'b 1000111000;
            10'b 1011000000 :   byte_offset = 10'b 1000111000;
            10'b 1011000001 :   byte_offset = 10'b 1000111001;
            10'b 1011000010 :   byte_offset = 10'b 1000111001;
            10'b 1011000011 :   byte_offset = 10'b 1000111010;
            10'b 1011000100 :   byte_offset = 10'b 1000111011;
            10'b 1011000101 :   byte_offset = 10'b 1000111011;
            10'b 1011000110 :   byte_offset = 10'b 1000111100;
            10'b 1011000111 :   byte_offset = 10'b 1000111100;
            10'b 1011001000 :   byte_offset = 10'b 1000111101;
            10'b 1011001001 :   byte_offset = 10'b 1000111101;
            10'b 1011001010 :   byte_offset = 10'b 1000111110;
            10'b 1011001011 :   byte_offset = 10'b 1000111111;
            10'b 1011001100 :   byte_offset = 10'b 1000111111;
            10'b 1011001101 :   byte_offset = 10'b 1001000000;
            10'b 1011001110 :   byte_offset = 10'b 1001000000;
            10'b 1011001111 :   byte_offset = 10'b 1001000001;
            10'b 1011010000 :   byte_offset = 10'b 1001000001;
            10'b 1011010001 :   byte_offset = 10'b 1001000010;
            10'b 1011010010 :   byte_offset = 10'b 1001000011;
            10'b 1011010011 :   byte_offset = 10'b 1001000011;
            10'b 1011010100 :   byte_offset = 10'b 1001000100;
            10'b 1011010101 :   byte_offset = 10'b 1001000100;
            10'b 1011010110 :   byte_offset = 10'b 1001000101;
            10'b 1011010111 :   byte_offset = 10'b 1001000101;
            10'b 1011011000 :   byte_offset = 10'b 1001010010;
            10'b 1011011001 :   byte_offset = 10'b 1001010011;
            10'b 1011011010 :   byte_offset = 10'b 1001010011;
            10'b 1011011011 :   byte_offset = 10'b 1001010100;
            10'b 1011011100 :   byte_offset = 10'b 1001010100;
            10'b 1011011101 :   byte_offset = 10'b 1001010101;
            10'b 1011011110 :   byte_offset = 10'b 1001010101;
            10'b 1011011111 :   byte_offset = 10'b 1001010110;
            10'b 1011100000 :   byte_offset = 10'b 1001010111;
            10'b 1011100001 :   byte_offset = 10'b 1001010111;
            10'b 1011100010 :   byte_offset = 10'b 1001011000;
            10'b 1011100011 :   byte_offset = 10'b 1001011000;
            10'b 1011100100 :   byte_offset = 10'b 1001011001;
            10'b 1011100101 :   byte_offset = 10'b 1001011001;
            10'b 1011100110 :   byte_offset = 10'b 1001011010;
            10'b 1011100111 :   byte_offset = 10'b 1001011011;
            10'b 1011101000 :   byte_offset = 10'b 1001011011;
            10'b 1011101001 :   byte_offset = 10'b 1001011100;
            10'b 1011101010 :   byte_offset = 10'b 1001011100;
            10'b 1011101011 :   byte_offset = 10'b 1001011101;
            10'b 1011101100 :   byte_offset = 10'b 1001011101;
            10'b 1011101101 :   byte_offset = 10'b 1001011110;
            10'b 1011101110 :   byte_offset = 10'b 1001011111;
            10'b 1011101111 :   byte_offset = 10'b 1001011111;
            10'b 1011110000 :   byte_offset = 10'b 1001100000;
            10'b 1011110001 :   byte_offset = 10'b 1001100000;
            10'b 1011110010 :   byte_offset = 10'b 1001100001;
            10'b 1011110011 :   byte_offset = 10'b 1001100001;
            10'b 1011110100 :   byte_offset = 10'b 1001010010;
            10'b 1011110101 :   byte_offset = 10'b 1001010011;
            10'b 1011110110 :   byte_offset = 10'b 1001010011;
            10'b 1011110111 :   byte_offset = 10'b 1001010100;
            10'b 1011111000 :   byte_offset = 10'b 1001010100;
            10'b 1011111001 :   byte_offset = 10'b 1001010101;
            10'b 1011111010 :   byte_offset = 10'b 1001010101;
            10'b 1011111011 :   byte_offset = 10'b 1001010110;
            10'b 1011111100 :   byte_offset = 10'b 1001010111;
            10'b 1011111101 :   byte_offset = 10'b 1001010111;
            10'b 1011111110 :   byte_offset = 10'b 1001011000;
            10'b 1011111111 :   byte_offset = 10'b 1001011000;
            10'b 1100000000 :   byte_offset = 10'b 1001011001;
            10'b 1100000001 :   byte_offset = 10'b 1001011001;
            10'b 1100000010 :   byte_offset = 10'b 1001011010;
            10'b 1100000011 :   byte_offset = 10'b 1001011011;
            10'b 1100000100 :   byte_offset = 10'b 1001011011;
            10'b 1100000101 :   byte_offset = 10'b 1001011100;
            10'b 1100000110 :   byte_offset = 10'b 1001011100;
            10'b 1100000111 :   byte_offset = 10'b 1001011101;
            10'b 1100001000 :   byte_offset = 10'b 1001011101;
            10'b 1100001001 :   byte_offset = 10'b 1001011110;
            10'b 1100001010 :   byte_offset = 10'b 1001011111;
            10'b 1100001011 :   byte_offset = 10'b 1001011111;
            10'b 1100001100 :   byte_offset = 10'b 1001100000;
            10'b 1100001101 :   byte_offset = 10'b 1001100000;
            10'b 1100001110 :   byte_offset = 10'b 1001100001;
            10'b 1100001111 :   byte_offset = 10'b 1001100001;
            default:            byte_offset = 10'b 0000000000;      

        endcase
    end
      assign address_offset = byte_offset;                      // add <<2 in case the bram is connected to PS instead of being an internal BRAM
endmodule