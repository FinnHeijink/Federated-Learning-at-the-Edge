module BRAM_sim_internal (
    input  logic [10:0] address,
    output logic [7:0]  data_send,
    input logic clk,
    input logic reset
);
    logic [7:0] data;
    
    always_ff @(posedge clk)
    if (reset)
    data_send <= 8'd0;
    else
    data_send <= data;





always_comb begin
    case (address)
        11'h000: data = 8'd0;
        11'h001: data = 8'd1;
        11'h002: data = 8'd2;
        11'h003: data = 8'd3;
        11'h004: data = 8'd4;
        11'h005: data = 8'd5;
        11'h006: data = 8'd6;
        11'h007: data = 8'd7;
        11'h008: data = 8'd8;
        11'h009: data = 8'd9;
        11'h00A: data = 8'd10;
        11'h00B: data = 8'd11;
        11'h00C: data = 8'd12;
        11'h00D: data = 8'd13;
        11'h00E: data = 8'd14;
        11'h00F: data = 8'd15;
        11'h010: data = 8'd16;
        11'h011: data = 8'd17;
        11'h012: data = 8'd18;
        11'h013: data = 8'd19;
        11'h014: data = 8'd20;
        11'h015: data = 8'd21;
        11'h016: data = 8'd22;
        11'h017: data = 8'd23;
        11'h018: data = 8'd24;
        11'h019: data = 8'd25;
        11'h01A: data = 8'd26;
        11'h01B: data = 8'd27;
        11'h01C: data = 8'd28;
        11'h01D: data = 8'd29;
        11'h01E: data = 8'd30;
        11'h01F: data = 8'd31;
        11'h020: data = 8'd32;
        11'h021: data = 8'd33;
        11'h022: data = 8'd34;
        11'h023: data = 8'd35;
        11'h024: data = 8'd36;
        11'h025: data = 8'd37;
        11'h026: data = 8'd38;
        11'h027: data = 8'd39;
        11'h028: data = 8'd40;
        11'h029: data = 8'd41;
        11'h02A: data = 8'd42;
        11'h02B: data = 8'd43;
        11'h02C: data = 8'd44;
        11'h02D: data = 8'd45;
        11'h02E: data = 8'd46;
        11'h02F: data = 8'd47;
        11'h030: data = 8'd48;
        11'h031: data = 8'd49;
        11'h032: data = 8'd50;
        11'h033: data = 8'd51;
        11'h034: data = 8'd52;
        11'h035: data = 8'd53;
        11'h036: data = 8'd54;
        11'h037: data = 8'd55;
        11'h038: data = 8'd56;
        11'h039: data = 8'd57;
        11'h03A: data = 8'd58;
        11'h03B: data = 8'd59;
        11'h03C: data = 8'd60;
        11'h03D: data = 8'd61;
        11'h03E: data = 8'd62;
        11'h03F: data = 8'd63;
        11'h040: data = 8'd64;
        11'h041: data = 8'd65;
        11'h042: data = 8'd66;
        11'h043: data = 8'd67;
        11'h044: data = 8'd68;
        11'h045: data = 8'd69;
        11'h046: data = 8'd70;
        11'h047: data = 8'd71;
        11'h048: data = 8'd72;
        11'h049: data = 8'd73;
        11'h04A: data = 8'd74;
        11'h04B: data = 8'd75;
        11'h04C: data = 8'd76;
        11'h04D: data = 8'd77;
        11'h04E: data = 8'd78;
        11'h04F: data = 8'd79;
        11'h050: data = 8'd80;
        11'h051: data = 8'd81;
        11'h052: data = 8'd82;
        11'h053: data = 8'd83;
        11'h054: data = 8'd84;
        11'h055: data = 8'd85;
        11'h056: data = 8'd86;
        11'h057: data = 8'd87;
        11'h058: data = 8'd88;
        11'h059: data = 8'd89;
        11'h05A: data = 8'd90;
        11'h05B: data = 8'd91;
        11'h05C: data = 8'd92;
        11'h05D: data = 8'd93;
        11'h05E: data = 8'd94;
        11'h05F: data = 8'd95;
        11'h060: data = 8'd96;
        11'h061: data = 8'd97;
        11'h062: data = 8'd98;
        11'h063: data = 8'd99;
        11'h064: data = 8'd100;
        11'h065: data = 8'd101;
        11'h066: data = 8'd102;
        11'h067: data = 8'd103;
        11'h068: data = 8'd104;
        11'h069: data = 8'd105;
        11'h06A: data = 8'd106;
        11'h06B: data = 8'd107;
        11'h06C: data = 8'd108;
        11'h06D: data = 8'd109;
        11'h06E: data = 8'd110;
        11'h06F: data = 8'd111;
        11'h070: data = 8'd112;
        11'h071: data = 8'd113;
        11'h072: data = 8'd114;
        11'h073: data = 8'd115;
        11'h074: data = 8'd116;
        11'h075: data = 8'd117;
        11'h076: data = 8'd118;
        11'h077: data = 8'd119;
        11'h078: data = 8'd120;
        11'h079: data = 8'd121;
        11'h07A: data = 8'd122;
        11'h07B: data = 8'd123;
        11'h07C: data = 8'd124;
        11'h07D: data = 8'd125;
        11'h07E: data = 8'd126;
        11'h07F: data = 8'd127;
        11'h080: data = 8'd128;
        11'h081: data = 8'd129;
        11'h082: data = 8'd130;
        11'h083: data = 8'd131;
        11'h084: data = 8'd132;
        11'h085: data = 8'd133;
        11'h086: data = 8'd134;
        11'h087: data = 8'd135;
        11'h088: data = 8'd136;
        11'h089: data = 8'd137;
        11'h08A: data = 8'd138;
        11'h08B: data = 8'd139;
        11'h08C: data = 8'd140;
        11'h08D: data = 8'd141;
        11'h08E: data = 8'd142;
        11'h08F: data = 8'd143;
        11'h090: data = 8'd144;
        11'h091: data = 8'd145;
        11'h092: data = 8'd146;
        11'h093: data = 8'd147;
        11'h094: data = 8'd148;
        11'h095: data = 8'd149;
        11'h096: data = 8'd150;
        11'h097: data = 8'd151;
        11'h098: data = 8'd152;
        11'h099: data = 8'd153;
        11'h09A: data = 8'd154;
        11'h09B: data = 8'd155;
        11'h09C: data = 8'd156;
        11'h09D: data = 8'd157;
        11'h09E: data = 8'd158;
        11'h09F: data = 8'd159;
        11'h0A0: data = 8'd160;
        11'h0A1: data = 8'd161;
        11'h0A2: data = 8'd162;
        11'h0A3: data = 8'd163;
        11'h0A4: data = 8'd164;
        11'h0A5: data = 8'd165;
        11'h0A6: data = 8'd166;
        11'h0A7: data = 8'd167;
        11'h0A8: data = 8'd168;
        11'h0A9: data = 8'd169;
        11'h0AA: data = 8'd170;
        11'h0AB: data = 8'd171;
        11'h0AC: data = 8'd172;
        11'h0AD: data = 8'd173;
        11'h0AE: data = 8'd174;
        11'h0AF: data = 8'd175;
        11'h0B0: data = 8'd176;
        11'h0B1: data = 8'd177;
        11'h0B2: data = 8'd178;
        11'h0B3: data = 8'd179;
        11'h0B4: data = 8'd180;
        11'h0B5: data = 8'd181;
        11'h0B6: data = 8'd182;
        11'h0B7: data = 8'd183;
        11'h0B8: data = 8'd184;
        11'h0B9: data = 8'd185;
        11'h0BA: data = 8'd186;
        11'h0BB: data = 8'd187;
        11'h0BC: data = 8'd188;
        11'h0BD: data = 8'd189;
        11'h0BE: data = 8'd190;
        11'h0BF: data = 8'd191;
        11'h0C0: data = 8'd192;
        11'h0C1: data = 8'd193;
        11'h0C2: data = 8'd194;
        11'h0C3: data = 8'd195;
        11'h0C4: data = 8'd196;
        11'h0C5: data = 8'd197;
        11'h0C6: data = 8'd198;
        11'h0C7: data = 8'd199;
        11'h0C8: data = 8'd200;
        11'h0C9: data = 8'd201;
        11'h0CA: data = 8'd202;
        11'h0CB: data = 8'd203;
        11'h0CC: data = 8'd204;
        11'h0CD: data = 8'd205;
        11'h0CE: data = 8'd206;
        11'h0CF: data = 8'd207;
        11'h0D0: data = 8'd208;
        11'h0D1: data = 8'd209;
        11'h0D2: data = 8'd210;
        11'h0D3: data = 8'd211;
        11'h0D4: data = 8'd212;
        11'h0D5: data = 8'd213;
        11'h0D6: data = 8'd214;
        11'h0D7: data = 8'd215;
        11'h0D8: data = 8'd216;
        11'h0D9: data = 8'd217;
        11'h0DA: data = 8'd218;
        11'h0DB: data = 8'd219;
        11'h0DC: data = 8'd220;
        11'h0DD: data = 8'd221;
        11'h0DE: data = 8'd222;
        11'h0DF: data = 8'd223;
        11'h0E0: data = 8'd224;
        11'h0E1: data = 8'd225;
        11'h0E2: data = 8'd226;
        11'h0E3: data = 8'd227;
        11'h0E4: data = 8'd228;
        11'h0E5: data = 8'd229;
        11'h0E6: data = 8'd230;
        11'h0E7: data = 8'd231;
        11'h0E8: data = 8'd232;
        11'h0E9: data = 8'd233;
        11'h0EA: data = 8'd234;
        11'h0EB: data = 8'd235;
        11'h0EC: data = 8'd236;
        11'h0ED: data = 8'd237;
        11'h0EE: data = 8'd238;
        11'h0EF: data = 8'd239;
        11'h0F0: data = 8'd240;
        11'h0F1: data = 8'd241;
        11'h0F2: data = 8'd242;
        11'h0F3: data = 8'd243;
        11'h0F4: data = 8'd244;
        11'h0F5: data = 8'd245;
        11'h0F6: data = 8'd246;
        11'h0F7: data = 8'd247;
        11'h0F8: data = 8'd248;
        11'h0F9: data = 8'd249;
        11'h0FA: data = 8'd250;
        11'h0FB: data = 8'd251;
        11'h0FC: data = 8'd252;
        11'h0FD: data = 8'd253;
        11'h0FE: data = 8'd254;
        11'h0FF: data = 8'd255;
        11'h100: data = 8'd256;
        11'h101: data = 8'd257;
        11'h102: data = 8'd258;
        11'h103: data = 8'd259;
        11'h104: data = 8'd260;
        11'h105: data = 8'd261;
        11'h106: data = 8'd262;
        11'h107: data = 8'd263;
        11'h108: data = 8'd264;
        11'h109: data = 8'd265;
        11'h10A: data = 8'd266;
        11'h10B: data = 8'd267;
        11'h10C: data = 8'd268;
        11'h10D: data = 8'd269;
        11'h10E: data = 8'd270;
        11'h10F: data = 8'd271;
        11'h110: data = 8'd272;
        11'h111: data = 8'd273;
        11'h112: data = 8'd274;
        11'h113: data = 8'd275;
        11'h114: data = 8'd276;
        11'h115: data = 8'd277;
        11'h116: data = 8'd278;
        11'h117: data = 8'd279;
        11'h118: data = 8'd280;
        11'h119: data = 8'd281;
        11'h11A: data = 8'd282;
        11'h11B: data = 8'd283;
        11'h11C: data = 8'd284;
        11'h11D: data = 8'd285;
        11'h11E: data = 8'd286;
        11'h11F: data = 8'd287;
        11'h120: data = 8'd288;
        11'h121: data = 8'd289;
        11'h122: data = 8'd290;
        11'h123: data = 8'd291;
        11'h124: data = 8'd292;
        11'h125: data = 8'd293;
        11'h126: data = 8'd294;
        11'h127: data = 8'd295;
        11'h128: data = 8'd296;
        11'h129: data = 8'd297;
        11'h12A: data = 8'd298;
        11'h12B: data = 8'd299;
        11'h12C: data = 8'd300;
        11'h12D: data = 8'd301;
        11'h12E: data = 8'd302;
        11'h12F: data = 8'd303;
        11'h130: data = 8'd304;
        11'h131: data = 8'd305;
        11'h132: data = 8'd306;
        11'h133: data = 8'd307;
        11'h134: data = 8'd308;
        11'h135: data = 8'd309;
        11'h136: data = 8'd310;
        11'h137: data = 8'd311;
        11'h138: data = 8'd312;
        11'h139: data = 8'd313;
        11'h13A: data = 8'd314;
        11'h13B: data = 8'd315;
        11'h13C: data = 8'd316;
        11'h13D: data = 8'd317;
        11'h13E: data = 8'd318;
        11'h13F: data = 8'd319;
        11'h140: data = 8'd320;
        11'h141: data = 8'd321;
        11'h142: data = 8'd322;
        11'h143: data = 8'd323;
        11'h144: data = 8'd324;
        11'h145: data = 8'd325;
        11'h146: data = 8'd326;
        11'h147: data = 8'd327;
        11'h148: data = 8'd328;
        11'h149: data = 8'd329;
        11'h14A: data = 8'd330;
        11'h14B: data = 8'd331;
        11'h14C: data = 8'd332;
        11'h14D: data = 8'd333;
        11'h14E: data = 8'd334;
        11'h14F: data = 8'd335;
        11'h150: data = 8'd336;
        11'h151: data = 8'd337;
        11'h152: data = 8'd338;
        11'h153: data = 8'd339;
        11'h154: data = 8'd340;
        11'h155: data = 8'd341;
        11'h156: data = 8'd342;
        11'h157: data = 8'd343;
        11'h158: data = 8'd344;
        11'h159: data = 8'd345;
        11'h15A: data = 8'd346;
        11'h15B: data = 8'd347;
        11'h15C: data = 8'd348;
        11'h15D: data = 8'd349;
        11'h15E: data = 8'd350;
        11'h15F: data = 8'd351;
        11'h160: data = 8'd352;
        11'h161: data = 8'd353;
        11'h162: data = 8'd354;
        11'h163: data = 8'd355;
        11'h164: data = 8'd356;
        11'h165: data = 8'd357;
        11'h166: data = 8'd358;
        11'h167: data = 8'd359;
        11'h168: data = 8'd360;
        11'h169: data = 8'd361;
        11'h16A: data = 8'd362;
        11'h16B: data = 8'd363;
        11'h16C: data = 8'd364;
        11'h16D: data = 8'd365;
        11'h16E: data = 8'd366;
        11'h16F: data = 8'd367;
        11'h170: data = 8'd368;
        11'h171: data = 8'd369;
        11'h172: data = 8'd370;
        11'h173: data = 8'd371;
        11'h174: data = 8'd372;
        11'h175: data = 8'd373;
        11'h176: data = 8'd374;
        11'h177: data = 8'd375;
        11'h178: data = 8'd376;
        11'h179: data = 8'd377;
        11'h17A: data = 8'd378;
        11'h17B: data = 8'd379;
        11'h17C: data = 8'd380;
        11'h17D: data = 8'd381;
        11'h17E: data = 8'd382;
        11'h17F: data = 8'd383;
        11'h180: data = 8'd384;
        11'h181: data = 8'd385;
        11'h182: data = 8'd386;
        11'h183: data = 8'd387;
        11'h184: data = 8'd388;
        11'h185: data = 8'd389;
        11'h186: data = 8'd390;
        11'h187: data = 8'd391;
        11'h188: data = 8'd392;
        11'h189: data = 8'd393;
        11'h18A: data = 8'd394;
        11'h18B: data = 8'd395;
        11'h18C: data = 8'd396;
        11'h18D: data = 8'd397;
        11'h18E: data = 8'd398;
        11'h18F: data = 8'd399;
        11'h190: data = 8'd400;
        11'h191: data = 8'd401;
        11'h192: data = 8'd402;
        11'h193: data = 8'd403;
        11'h194: data = 8'd404;
        11'h195: data = 8'd405;
        11'h196: data = 8'd406;
        11'h197: data = 8'd407;
        11'h198: data = 8'd408;
        11'h199: data = 8'd409;
        11'h19A: data = 8'd410;
        11'h19B: data = 8'd411;
        11'h19C: data = 8'd412;
        11'h19D: data = 8'd413;
        11'h19E: data = 8'd414;
        11'h19F: data = 8'd415;
        11'h1A0: data = 8'd416;
        11'h1A1: data = 8'd417;
        11'h1A2: data = 8'd418;
        11'h1A3: data = 8'd419;
        11'h1A4: data = 8'd420;
        11'h1A5: data = 8'd421;
        11'h1A6: data = 8'd422;
        11'h1A7: data = 8'd423;
        11'h1A8: data = 8'd424;
        11'h1A9: data = 8'd425;
        11'h1AA: data = 8'd426;
        11'h1AB: data = 8'd427;
        11'h1AC: data = 8'd428;
        11'h1AD: data = 8'd429;
        11'h1AE: data = 8'd430;
        11'h1AF: data = 8'd431;
        11'h1B0: data = 8'd432;
        11'h1B1: data = 8'd433;
        11'h1B2: data = 8'd434;
        11'h1B3: data = 8'd435;
        11'h1B4: data = 8'd436;
        11'h1B5: data = 8'd437;
        11'h1B6: data = 8'd438;
        11'h1B7: data = 8'd439;
        11'h1B8: data = 8'd440;
        11'h1B9: data = 8'd441;
        11'h1BA: data = 8'd442;
        11'h1BB: data = 8'd443;
        11'h1BC: data = 8'd444;
        11'h1BD: data = 8'd445;
        11'h1BE: data = 8'd446;
        11'h1BF: data = 8'd447;
        11'h1C0: data = 8'd448;
        11'h1C1: data = 8'd449;
        11'h1C2: data = 8'd450;
        11'h1C3: data = 8'd451;
        11'h1C4: data = 8'd452;
        11'h1C5: data = 8'd453;
        11'h1C6: data = 8'd454;
        11'h1C7: data = 8'd455;
        11'h1C8: data = 8'd456;
        11'h1C9: data = 8'd457;
        11'h1CA: data = 8'd458;
        11'h1CB: data = 8'd459;
        11'h1CC: data = 8'd460;
        11'h1CD: data = 8'd461;
        11'h1CE: data = 8'd462;
        11'h1CF: data = 8'd463;
        11'h1D0: data = 8'd464;
        11'h1D1: data = 8'd465;
        11'h1D2: data = 8'd466;
        11'h1D3: data = 8'd467;
        11'h1D4: data = 8'd468;
        11'h1D5: data = 8'd469;
        11'h1D6: data = 8'd470;
        11'h1D7: data = 8'd471;
        11'h1D8: data = 8'd472;
        11'h1D9: data = 8'd473;
        11'h1DA: data = 8'd474;
        11'h1DB: data = 8'd475;
        11'h1DC: data = 8'd476;
        11'h1DD: data = 8'd477;
        11'h1DE: data = 8'd478;
        11'h1DF: data = 8'd479;
        11'h1E0: data = 8'd480;
        11'h1E1: data = 8'd481;
        11'h1E2: data = 8'd482;
        11'h1E3: data = 8'd483;
        11'h1E4: data = 8'd484;
        11'h1E5: data = 8'd485;
        11'h1E6: data = 8'd486;
        11'h1E7: data = 8'd487;
        11'h1E8: data = 8'd488;
        11'h1E9: data = 8'd489;
        11'h1EA: data = 8'd490;
        11'h1EB: data = 8'd491;
        11'h1EC: data = 8'd492;
        11'h1ED: data = 8'd493;
        11'h1EE: data = 8'd494;
        11'h1EF: data = 8'd495;
        11'h1F0: data = 8'd496;
        11'h1F1: data = 8'd497;
        11'h1F2: data = 8'd498;
        11'h1F3: data = 8'd499;
        11'h1F4: data = 8'd500;
        11'h1F5: data = 8'd501;
        11'h1F6: data = 8'd502;
        11'h1F7: data = 8'd503;
        11'h1F8: data = 8'd504;
        11'h1F9: data = 8'd505;
        11'h1FA: data = 8'd506;
        11'h1FB: data = 8'd507;
        11'h1FC: data = 8'd508;
        11'h1FD: data = 8'd509;
        11'h1FE: data = 8'd510;
        11'h1FF: data = 8'd511;
        11'h200: data = 8'd512;
        11'h201: data = 8'd513;
        11'h202: data = 8'd514;
        11'h203: data = 8'd515;
        11'h204: data = 8'd516;
        11'h205: data = 8'd517;
        11'h206: data = 8'd518;
        11'h207: data = 8'd519;
        11'h208: data = 8'd520;
        11'h209: data = 8'd521;
        11'h20A: data = 8'd522;
        11'h20B: data = 8'd523;
        11'h20C: data = 8'd524;
        11'h20D: data = 8'd525;
        11'h20E: data = 8'd526;
        11'h20F: data = 8'd527;
        11'h210: data = 8'd528;
        11'h211: data = 8'd529;
        11'h212: data = 8'd530;
        11'h213: data = 8'd531;
        11'h214: data = 8'd532;
        11'h215: data = 8'd533;
        11'h216: data = 8'd534;
        11'h217: data = 8'd535;
        11'h218: data = 8'd536;
        11'h219: data = 8'd537;
        11'h21A: data = 8'd538;
        11'h21B: data = 8'd539;
        11'h21C: data = 8'd540;
        11'h21D: data = 8'd541;
        11'h21E: data = 8'd542;
        11'h21F: data = 8'd543;
        11'h220: data = 8'd544;
        11'h221: data = 8'd545;
        11'h222: data = 8'd546;
        11'h223: data = 8'd547;
        11'h224: data = 8'd548;
        11'h225: data = 8'd549;
        11'h226: data = 8'd550;
        11'h227: data = 8'd551;
        11'h228: data = 8'd552;
        11'h229: data = 8'd553;
        11'h22A: data = 8'd554;
        11'h22B: data = 8'd555;
        11'h22C: data = 8'd556;
        11'h22D: data = 8'd557;
        11'h22E: data = 8'd558;
        11'h22F: data = 8'd559;
        11'h230: data = 8'd560;
        11'h231: data = 8'd561;
        11'h232: data = 8'd562;
        11'h233: data = 8'd563;
        11'h234: data = 8'd564;
        11'h235: data = 8'd565;
        11'h236: data = 8'd566;
        11'h237: data = 8'd567;
        11'h238: data = 8'd568;
        11'h239: data = 8'd569;
        11'h23A: data = 8'd570;
        11'h23B: data = 8'd571;
        11'h23C: data = 8'd572;
        11'h23D: data = 8'd573;
        11'h23E: data = 8'd574;
        11'h23F: data = 8'd575;
        11'h240: data = 8'd576;
        11'h241: data = 8'd577;
        11'h242: data = 8'd578;
        11'h243: data = 8'd579;
        11'h244: data = 8'd580;
        11'h245: data = 8'd581;
        11'h246: data = 8'd582;
        11'h247: data = 8'd583;
        11'h248: data = 8'd584;
        11'h249: data = 8'd585;
        11'h24A: data = 8'd586;
        11'h24B: data = 8'd587;
        11'h24C: data = 8'd588;
        11'h24D: data = 8'd589;
        11'h24E: data = 8'd590;
        11'h24F: data = 8'd591;
        11'h250: data = 8'd592;
        11'h251: data = 8'd593;
        11'h252: data = 8'd594;
        11'h253: data = 8'd595;
        11'h254: data = 8'd596;
        11'h255: data = 8'd597;
        11'h256: data = 8'd598;
        11'h257: data = 8'd599;
        11'h258: data = 8'd600;
        11'h259: data = 8'd601;
        11'h25A: data = 8'd602;
        11'h25B: data = 8'd603;
        11'h25C: data = 8'd604;
        11'h25D: data = 8'd605;
        11'h25E: data = 8'd606;
        11'h25F: data = 8'd607;
        11'h260: data = 8'd608;
        11'h261: data = 8'd609;
        11'h262: data = 8'd610;
        11'h263: data = 8'd611;
        11'h264: data = 8'd612;
        11'h265: data = 8'd613;
        11'h266: data = 8'd614;
        11'h267: data = 8'd615;
        11'h268: data = 8'd616;
        11'h269: data = 8'd617;
        11'h26A: data = 8'd618;
        11'h26B: data = 8'd619;
        11'h26C: data = 8'd620;
        11'h26D: data = 8'd621;
        11'h26E: data = 8'd622;
        11'h26F: data = 8'd623;
        11'h270: data = 8'd624;
        11'h271: data = 8'd625;
        11'h272: data = 8'd626;
        11'h273: data = 8'd627;
        11'h274: data = 8'd628;
        11'h275: data = 8'd629;
        11'h276: data = 8'd630;
        11'h277: data = 8'd631;
        11'h278: data = 8'd632;
        11'h279: data = 8'd633;
        11'h27A: data = 8'd634;
        11'h27B: data = 8'd635;
        11'h27C: data = 8'd636;
        11'h27D: data = 8'd637;
        11'h27E: data = 8'd638;
        11'h27F: data = 8'd639;
        11'h280: data = 8'd640;
        11'h281: data = 8'd641;
        11'h282: data = 8'd642;
        11'h283: data = 8'd643;
        11'h284: data = 8'd644;
        11'h285: data = 8'd645;
        11'h286: data = 8'd646;
        11'h287: data = 8'd647;
        11'h288: data = 8'd648;
        11'h289: data = 8'd649;
        11'h28A: data = 8'd650;
        11'h28B: data = 8'd651;
        11'h28C: data = 8'd652;
        11'h28D: data = 8'd653;
        11'h28E: data = 8'd654;
        11'h28F: data = 8'd655;
        11'h290: data = 8'd656;
        11'h291: data = 8'd657;
        11'h292: data = 8'd658;
        11'h293: data = 8'd659;
        11'h294: data = 8'd660;
        11'h295: data = 8'd661;
        11'h296: data = 8'd662;
        11'h297: data = 8'd663;
        11'h298: data = 8'd664;
        11'h299: data = 8'd665;
        11'h29A: data = 8'd666;
        11'h29B: data = 8'd667;
        11'h29C: data = 8'd668;
        11'h29D: data = 8'd669;
        11'h29E: data = 8'd670;
        11'h29F: data = 8'd671;
        11'h2A0: data = 8'd672;
        11'h2A1: data = 8'd673;
        11'h2A2: data = 8'd674;
        11'h2A3: data = 8'd675;
        11'h2A4: data = 8'd676;
        11'h2A5: data = 8'd677;
        11'h2A6: data = 8'd678;
        11'h2A7: data = 8'd679;
        11'h2A8: data = 8'd680;
        11'h2A9: data = 8'd681;
        11'h2AA: data = 8'd682;
        11'h2AB: data = 8'd683;
        11'h2AC: data = 8'd684;
        11'h2AD: data = 8'd685;
        11'h2AE: data = 8'd686;
        11'h2AF: data = 8'd687;
        11'h2B0: data = 8'd688;
        11'h2B1: data = 8'd689;
        11'h2B2: data = 8'd690;
        11'h2B3: data = 8'd691;
        11'h2B4: data = 8'd692;
        11'h2B5: data = 8'd693;
        11'h2B6: data = 8'd694;
        11'h2B7: data = 8'd695;
        11'h2B8: data = 8'd696;
        11'h2B9: data = 8'd697;
        11'h2BA: data = 8'd698;
        11'h2BB: data = 8'd699;
        11'h2BC: data = 8'd700;
        11'h2BD: data = 8'd701;
        11'h2BE: data = 8'd702;
        11'h2BF: data = 8'd703;
        11'h2C0: data = 8'd704;
        11'h2C1: data = 8'd705;
        11'h2C2: data = 8'd706;
        11'h2C3: data = 8'd707;
        11'h2C4: data = 8'd708;
        11'h2C5: data = 8'd709;
        11'h2C6: data = 8'd710;
        11'h2C7: data = 8'd711;
        11'h2C8: data = 8'd712;
        11'h2C9: data = 8'd713;
        11'h2CA: data = 8'd714;
        11'h2CB: data = 8'd715;
        11'h2CC: data = 8'd716;
        11'h2CD: data = 8'd717;
        11'h2CE: data = 8'd718;
        11'h2CF: data = 8'd719;
        11'h2D0: data = 8'd720;
        11'h2D1: data = 8'd721;
        11'h2D2: data = 8'd722;
        11'h2D3: data = 8'd723;
        11'h2D4: data = 8'd724;
        11'h2D5: data = 8'd725;
        11'h2D6: data = 8'd726;
        11'h2D7: data = 8'd727;
        11'h2D8: data = 8'd728;
        11'h2D9: data = 8'd729;
        11'h2DA: data = 8'd730;
        11'h2DB: data = 8'd731;
        11'h2DC: data = 8'd732;
        11'h2DD: data = 8'd733;
        11'h2DE: data = 8'd734;
        11'h2DF: data = 8'd735;
        11'h2E0: data = 8'd736;
        11'h2E1: data = 8'd737;
        11'h2E2: data = 8'd738;
        11'h2E3: data = 8'd739;
        11'h2E4: data = 8'd740;
        11'h2E5: data = 8'd741;
        11'h2E6: data = 8'd742;
        11'h2E7: data = 8'd743;
        11'h2E8: data = 8'd744;
        11'h2E9: data = 8'd745;
        11'h2EA: data = 8'd746;
        11'h2EB: data = 8'd747;
        11'h2EC: data = 8'd748;
        11'h2ED: data = 8'd749;
        11'h2EE: data = 8'd750;
        11'h2EF: data = 8'd751;
        11'h2F0: data = 8'd752;
        11'h2F1: data = 8'd753;
        11'h2F2: data = 8'd754;
        11'h2F3: data = 8'd755;
        11'h2F4: data = 8'd756;
        11'h2F5: data = 8'd757;
        11'h2F6: data = 8'd758;
        11'h2F7: data = 8'd759;
        11'h2F8: data = 8'd760;
        11'h2F9: data = 8'd761;
        11'h2FA: data = 8'd762;
        11'h2FB: data = 8'd763;
        11'h2FC: data = 8'd764;
        11'h2FD: data = 8'd765;
        11'h2FE: data = 8'd766;
        11'h2FF: data = 8'd767;
        11'h300: data = 8'd768;
        11'h301: data = 8'd769;
        11'h302: data = 8'd770;
        11'h303: data = 8'd771;
        11'h304: data = 8'd772;
        11'h305: data = 8'd773;
        11'h306: data = 8'd774;
        11'h307: data = 8'd775;
        11'h308: data = 8'd776;
        11'h309: data = 8'd777;
        11'h30A: data = 8'd778;
        11'h30B: data = 8'd779;
        11'h30C: data = 8'd780;
        11'h30D: data = 8'd781;
        11'h30E: data = 8'd782;
        11'h30F: data = 8'd783;
        11'h310: data = 8'd784;
        11'h311: data = 8'd785;
        11'h312: data = 8'd786;
        11'h313: data = 8'd787;
        11'h314: data = 8'd788;
        11'h315: data = 8'd789;
        11'h316: data = 8'd790;
        11'h317: data = 8'd791;
        11'h318: data = 8'd792;
        11'h319: data = 8'd793;
        11'h31A: data = 8'd794;
        11'h31B: data = 8'd795;
        11'h31C: data = 8'd796;
        11'h31D: data = 8'd797;
        11'h31E: data = 8'd798;
        11'h31F: data = 8'd799;
        11'h320: data = 8'd800;
        11'h321: data = 8'd801;
        11'h322: data = 8'd802;
        11'h323: data = 8'd803;
        11'h324: data = 8'd804;
        11'h325: data = 8'd805;
        11'h326: data = 8'd806;
        11'h327: data = 8'd807;
        11'h328: data = 8'd808;
        11'h329: data = 8'd809;
        11'h32A: data = 8'd810;
        11'h32B: data = 8'd811;
        11'h32C: data = 8'd812;
        11'h32D: data = 8'd813;
        11'h32E: data = 8'd814;
        11'h32F: data = 8'd815;
        11'h330: data = 8'd816;
        11'h331: data = 8'd817;
        11'h332: data = 8'd818;
        11'h333: data = 8'd819;
        11'h334: data = 8'd820;
        11'h335: data = 8'd821;
        11'h336: data = 8'd822;
        11'h337: data = 8'd823;
        11'h338: data = 8'd824;
        11'h339: data = 8'd825;
        11'h33A: data = 8'd826;
        11'h33B: data = 8'd827;
        11'h33C: data = 8'd828;
        11'h33D: data = 8'd829;
        11'h33E: data = 8'd830;
        11'h33F: data = 8'd831;
        11'h340: data = 8'd832;
        11'h341: data = 8'd833;
        11'h342: data = 8'd834;
        11'h343: data = 8'd835;
        11'h344: data = 8'd836;
        11'h345: data = 8'd837;
        11'h346: data = 8'd838;
        11'h347: data = 8'd839;
        11'h348: data = 8'd840;
        11'h349: data = 8'd841;
        11'h34A: data = 8'd842;
        11'h34B: data = 8'd843;
        11'h34C: data = 8'd844;
        11'h34D: data = 8'd845;
        11'h34E: data = 8'd846;
        11'h34F: data = 8'd847;
        11'h350: data = 8'd848;
        11'h351: data = 8'd849;
        11'h352: data = 8'd850;
        11'h353: data = 8'd851;
        11'h354: data = 8'd852;
        11'h355: data = 8'd853;
        11'h356: data = 8'd854;
        11'h357: data = 8'd855;
        11'h358: data = 8'd856;
        11'h359: data = 8'd857;
        11'h35A: data = 8'd858;
        11'h35B: data = 8'd859;
        11'h35C: data = 8'd860;
        11'h35D: data = 8'd861;
        11'h35E: data = 8'd862;
        11'h35F: data = 8'd863;
        11'h360: data = 8'd864;
        11'h361: data = 8'd865;
        11'h362: data = 8'd866;
        11'h363: data = 8'd867;
        11'h364: data = 8'd868;
        11'h365: data = 8'd869;
        11'h366: data = 8'd870;
        11'h367: data = 8'd871;
        11'h368: data = 8'd872;
        11'h369: data = 8'd873;
        11'h36A: data = 8'd874;
        11'h36B: data = 8'd875;
        11'h36C: data = 8'd876;
        11'h36D: data = 8'd877;
        11'h36E: data = 8'd878;
        11'h36F: data = 8'd879;
        11'h370: data = 8'd880;
        11'h371: data = 8'd881;
        11'h372: data = 8'd882;
        11'h373: data = 8'd883;
        11'h374: data = 8'd884;
        11'h375: data = 8'd885;
        11'h376: data = 8'd886;
        11'h377: data = 8'd887;
        11'h378: data = 8'd888;
        11'h379: data = 8'd889;
        11'h37A: data = 8'd890;
        11'h37B: data = 8'd891;
        11'h37C: data = 8'd892;
        11'h37D: data = 8'd893;
        11'h37E: data = 8'd894;
        11'h37F: data = 8'd895;
        11'h380: data = 8'd896;
        11'h381: data = 8'd897;
        11'h382: data = 8'd898;
        11'h383: data = 8'd899;
        11'h384: data = 8'd900;
        11'h385: data = 8'd901;
        11'h386: data = 8'd902;
        11'h387: data = 8'd903;
        11'h388: data = 8'd904;
        11'h389: data = 8'd905;
        11'h38A: data = 8'd906;
        11'h38B: data = 8'd907;
        11'h38C: data = 8'd908;
        11'h38D: data = 8'd909;
        11'h38E: data = 8'd910;
        11'h38F: data = 8'd911;
        11'h390: data = 8'd912;
        11'h391: data = 8'd913;
        11'h392: data = 8'd914;
        11'h393: data = 8'd915;
        11'h394: data = 8'd916;
        11'h395: data = 8'd917;
        11'h396: data = 8'd918;
        11'h397: data = 8'd919;
        11'h398: data = 8'd920;
        11'h399: data = 8'd921;
        11'h39A: data = 8'd922;
        11'h39B: data = 8'd923;
        11'h39C: data = 8'd924;
        11'h39D: data = 8'd925;
        11'h39E: data = 8'd926;
        11'h39F: data = 8'd927;
        11'h3A0: data = 8'd928;
        11'h3A1: data = 8'd929;
        11'h3A2: data = 8'd930;
        11'h3A3: data = 8'd931;
        11'h3A4: data = 8'd932;
        11'h3A5: data = 8'd933;
        11'h3A6: data = 8'd934;
        11'h3A7: data = 8'd935;
        11'h3A8: data = 8'd936;
        11'h3A9: data = 8'd937;
        11'h3AA: data = 8'd938;
        11'h3AB: data = 8'd939;
        11'h3AC: data = 8'd940;
        11'h3AD: data = 8'd941;
        11'h3AE: data = 8'd942;
        11'h3AF: data = 8'd943;
        11'h3B0: data = 8'd944;
        11'h3B1: data = 8'd945;
        11'h3B2: data = 8'd946;
        11'h3B3: data = 8'd947;
        11'h3B4: data = 8'd948;
        11'h3B5: data = 8'd949;
        11'h3B6: data = 8'd950;
        11'h3B7: data = 8'd951;
        11'h3B8: data = 8'd952;
        11'h3B9: data = 8'd953;
        11'h3BA: data = 8'd954;
        11'h3BB: data = 8'd955;
        11'h3BC: data = 8'd956;
        11'h3BD: data = 8'd957;
        11'h3BE: data = 8'd958;
        11'h3BF: data = 8'd959;
        11'h3C0: data = 8'd960;
        11'h3C1: data = 8'd961;
        11'h3C2: data = 8'd962;
        11'h3C3: data = 8'd963;
        11'h3C4: data = 8'd964;
        11'h3C5: data = 8'd965;
        11'h3C6: data = 8'd966;
        11'h3C7: data = 8'd967;
        11'h3C8: data = 8'd968;
        11'h3C9: data = 8'd969;
        11'h3CA: data = 8'd970;
        11'h3CB: data = 8'd971;
        11'h3CC: data = 8'd972;
        11'h3CD: data = 8'd973;
        11'h3CE: data = 8'd974;
        11'h3CF: data = 8'd975;
        11'h3D0: data = 8'd976;
        11'h3D1: data = 8'd977;
        11'h3D2: data = 8'd978;
        11'h3D3: data = 8'd979;
        11'h3D4: data = 8'd980;
        11'h3D5: data = 8'd981;
        11'h3D6: data = 8'd982;
        11'h3D7: data = 8'd983;
        11'h3D8: data = 8'd984;
        11'h3D9: data = 8'd985;
        11'h3DA: data = 8'd986;
        11'h3DB: data = 8'd987;
        11'h3DC: data = 8'd988;
        11'h3DD: data = 8'd989;
        11'h3DE: data = 8'd990;
        11'h3DF: data = 8'd991;
        11'h3E0: data = 8'd992;
        11'h3E1: data = 8'd993;
        11'h3E2: data = 8'd994;
        11'h3E3: data = 8'd995;
        11'h3E4: data = 8'd996;
        11'h3E5: data = 8'd997;
        11'h3E6: data = 8'd998;
        11'h3E7: data = 8'd999;
        11'h3E8: data = 8'd1000;
        11'h3E9: data = 8'd1001;
        11'h3EA: data = 8'd1002;
        11'h3EB: data = 8'd1003;
        11'h3EC: data = 8'd1004;
        11'h3ED: data = 8'd1005;
        11'h3EE: data = 8'd1006;
        11'h3EF: data = 8'd1007;
        11'h3F0: data = 8'd1008;
        11'h3F1: data = 8'd1009;
        11'h3F2: data = 8'd1010;
        11'h3F3: data = 8'd1011;
        11'h3F4: data = 8'd1012;
        11'h3F5: data = 8'd1013;
        11'h3F6: data = 8'd1014;
        11'h3F7: data = 8'd1015;
        11'h3F8: data = 8'd1016;
        11'h3F9: data = 8'd1017;
        11'h3FA: data = 8'd1018;
        11'h3FB: data = 8'd1019;
        11'h3FC: data = 8'd1020;
        11'h3FD: data = 8'd1021;
        11'h3FE: data = 8'd1022;
        11'h3FF: data = 8'd1023;
        11'h400: data = 8'd1024;
        11'h401: data = 8'd1025;
        11'h402: data = 8'd1026;
        11'h403: data = 8'd1027;
        11'h404: data = 8'd1028;
        11'h405: data = 8'd1029;
        11'h406: data = 8'd1030;
        11'h407: data = 8'd1031;
        11'h408: data = 8'd1032;
        11'h409: data = 8'd1033;
        11'h40A: data = 8'd1034;
        11'h40B: data = 8'd1035;
        11'h40C: data = 8'd1036;
        11'h40D: data = 8'd1037;
        11'h40E: data = 8'd1038;
        11'h40F: data = 8'd1039;
        11'h410: data = 8'd1040;
        11'h411: data = 8'd1041;
        11'h412: data = 8'd1042;
        11'h413: data = 8'd1043;
        11'h414: data = 8'd1044;
        11'h415: data = 8'd1045;
        11'h416: data = 8'd1046;
        11'h417: data = 8'd1047;
        11'h418: data = 8'd1048;
        11'h419: data = 8'd1049;
        11'h41A: data = 8'd1050;
        11'h41B: data = 8'd1051;
        11'h41C: data = 8'd1052;
        11'h41D: data = 8'd1053;
        11'h41E: data = 8'd1054;
        11'h41F: data = 8'd1055;
        11'h420: data = 8'd1056;
        11'h421: data = 8'd1057;
        11'h422: data = 8'd1058;
        11'h423: data = 8'd1059;
        11'h424: data = 8'd1060;
        11'h425: data = 8'd1061;
        11'h426: data = 8'd1062;
        11'h427: data = 8'd1063;
        11'h428: data = 8'd1064;
        11'h429: data = 8'd1065;
        11'h42A: data = 8'd1066;
        11'h42B: data = 8'd1067;
        11'h42C: data = 8'd1068;
        11'h42D: data = 8'd1069;
        11'h42E: data = 8'd1070;
        11'h42F: data = 8'd1071;
        11'h430: data = 8'd1072;
        11'h431: data = 8'd1073;
        11'h432: data = 8'd1074;
        11'h433: data = 8'd1075;
        11'h434: data = 8'd1076;
        11'h435: data = 8'd1077;
        11'h436: data = 8'd1078;
        11'h437: data = 8'd1079;
        11'h438: data = 8'd1080;
        11'h439: data = 8'd1081;
        11'h43A: data = 8'd1082;
        11'h43B: data = 8'd1083;
        11'h43C: data = 8'd1084;
        11'h43D: data = 8'd1085;
        11'h43E: data = 8'd1086;
        11'h43F: data = 8'd1087;
        11'h440: data = 8'd1088;
        11'h441: data = 8'd1089;
        11'h442: data = 8'd1090;
        11'h443: data = 8'd1091;
        11'h444: data = 8'd1092;
        11'h445: data = 8'd1093;
        11'h446: data = 8'd1094;
        11'h447: data = 8'd1095;
        11'h448: data = 8'd1096;
        11'h449: data = 8'd1097;
        11'h44A: data = 8'd1098;
        11'h44B: data = 8'd1099;
        11'h44C: data = 8'd1100;
        11'h44D: data = 8'd1101;
        11'h44E: data = 8'd1102;
        11'h44F: data = 8'd1103;
        11'h450: data = 8'd1104;
        11'h451: data = 8'd1105;
        11'h452: data = 8'd1106;
        11'h453: data = 8'd1107;
        11'h454: data = 8'd1108;
        11'h455: data = 8'd1109;
        11'h456: data = 8'd1110;
        11'h457: data = 8'd1111;
        11'h458: data = 8'd1112;
        11'h459: data = 8'd1113;
        11'h45A: data = 8'd1114;
        11'h45B: data = 8'd1115;
        11'h45C: data = 8'd1116;
        11'h45D: data = 8'd1117;
        11'h45E: data = 8'd1118;
        11'h45F: data = 8'd1119;
        11'h460: data = 8'd1120;
        11'h461: data = 8'd1121;
        11'h462: data = 8'd1122;
        11'h463: data = 8'd1123;
        11'h464: data = 8'd1124;
        11'h465: data = 8'd1125;
        11'h466: data = 8'd1126;
        11'h467: data = 8'd1127;
        11'h468: data = 8'd1128;
        11'h469: data = 8'd1129;
        11'h46A: data = 8'd1130;
        11'h46B: data = 8'd1131;
        11'h46C: data = 8'd1132;
        11'h46D: data = 8'd1133;
        11'h46E: data = 8'd1134;
        11'h46F: data = 8'd1135;
        11'h470: data = 8'd1136;
        11'h471: data = 8'd1137;
        11'h472: data = 8'd1138;
        11'h473: data = 8'd1139;
        11'h474: data = 8'd1140;
        11'h475: data = 8'd1141;
        11'h476: data = 8'd1142;
        11'h477: data = 8'd1143;
        11'h478: data = 8'd1144;
        11'h479: data = 8'd1145;
        11'h47A: data = 8'd1146;
        11'h47B: data = 8'd1147;
        11'h47C: data = 8'd1148;
        11'h47D: data = 8'd1149;
        11'h47E: data = 8'd1150;
        11'h47F: data = 8'd1151;
        11'h480: data = 8'd1152;
        11'h481: data = 8'd1153;
        11'h482: data = 8'd1154;
        11'h483: data = 8'd1155;
        11'h484: data = 8'd1156;
        11'h485: data = 8'd1157;
        11'h486: data = 8'd1158;
        11'h487: data = 8'd1159;
        11'h488: data = 8'd1160;
        11'h489: data = 8'd1161;
        11'h48A: data = 8'd1162;
        11'h48B: data = 8'd1163;
        11'h48C: data = 8'd1164;
        11'h48D: data = 8'd1165;
        11'h48E: data = 8'd1166;
        11'h48F: data = 8'd1167;
        11'h490: data = 8'd1168;
        11'h491: data = 8'd1169;
        11'h492: data = 8'd1170;
        11'h493: data = 8'd1171;
        11'h494: data = 8'd1172;
        11'h495: data = 8'd1173;
        11'h496: data = 8'd1174;
        11'h497: data = 8'd1175;
        11'h498: data = 8'd1176;
        11'h499: data = 8'd1177;
        11'h49A: data = 8'd1178;
        11'h49B: data = 8'd1179;
        11'h49C: data = 8'd1180;
        11'h49D: data = 8'd1181;
        11'h49E: data = 8'd1182;
        11'h49F: data = 8'd1183;
        11'h4A0: data = 8'd1184;
        11'h4A1: data = 8'd1185;
        11'h4A2: data = 8'd1186;
        11'h4A3: data = 8'd1187;
        11'h4A4: data = 8'd1188;
        11'h4A5: data = 8'd1189;
        11'h4A6: data = 8'd1190;
        11'h4A7: data = 8'd1191;
        11'h4A8: data = 8'd1192;
        11'h4A9: data = 8'd1193;
        11'h4AA: data = 8'd1194;
        11'h4AB: data = 8'd1195;
        11'h4AC: data = 8'd1196;
        11'h4AD: data = 8'd1197;
        11'h4AE: data = 8'd1198;
        11'h4AF: data = 8'd1199;
        11'h4B0: data = 8'd1200;
        11'h4B1: data = 8'd1201;
        11'h4B2: data = 8'd1202;
        11'h4B3: data = 8'd1203;
        11'h4B4: data = 8'd1204;
        11'h4B5: data = 8'd1205;
        11'h4B6: data = 8'd1206;
        11'h4B7: data = 8'd1207;
        11'h4B8: data = 8'd1208;
        11'h4B9: data = 8'd1209;
        11'h4BA: data = 8'd1210;
        11'h4BB: data = 8'd1211;
        11'h4BC: data = 8'd1212;
        11'h4BD: data = 8'd1213;
        11'h4BE: data = 8'd1214;
        11'h4BF: data = 8'd1215;
        11'h4C0: data = 8'd1216;
        11'h4C1: data = 8'd1217;
        11'h4C2: data = 8'd1218;
        11'h4C3: data = 8'd1219;
        11'h4C4: data = 8'd1220;
        11'h4C5: data = 8'd1221;
        11'h4C6: data = 8'd1222;
        11'h4C7: data = 8'd1223;
        11'h4C8: data = 8'd1224;
        11'h4C9: data = 8'd1225;
        11'h4CA: data = 8'd1226;
        11'h4CB: data = 8'd1227;
        11'h4CC: data = 8'd1228;
        11'h4CD: data = 8'd1229;
        11'h4CE: data = 8'd1230;
        11'h4CF: data = 8'd1231;
        11'h4D0: data = 8'd1232;
        11'h4D1: data = 8'd1233;
        11'h4D2: data = 8'd1234;
        11'h4D3: data = 8'd1235;
        11'h4D4: data = 8'd1236;
        11'h4D5: data = 8'd1237;
        11'h4D6: data = 8'd1238;
        11'h4D7: data = 8'd1239;
        11'h4D8: data = 8'd1240;
        11'h4D9: data = 8'd1241;
        11'h4DA: data = 8'd1242;
        11'h4DB: data = 8'd1243;
        11'h4DC: data = 8'd1244;
        11'h4DD: data = 8'd1245;
        11'h4DE: data = 8'd1246;
        11'h4DF: data = 8'd1247;
        11'h4E0: data = 8'd1248;
        11'h4E1: data = 8'd1249;
        11'h4E2: data = 8'd1250;
        11'h4E3: data = 8'd1251;
        11'h4E4: data = 8'd1252;
        11'h4E5: data = 8'd1253;
        11'h4E6: data = 8'd1254;
        11'h4E7: data = 8'd1255;
        11'h4E8: data = 8'd1256;
        11'h4E9: data = 8'd1257;
        11'h4EA: data = 8'd1258;
        11'h4EB: data = 8'd1259;
        11'h4EC: data = 8'd1260;
        11'h4ED: data = 8'd1261;
        11'h4EE: data = 8'd1262;
        11'h4EF: data = 8'd1263;
        11'h4F0: data = 8'd1264;
        11'h4F1: data = 8'd1265;
        11'h4F2: data = 8'd1266;
        11'h4F3: data = 8'd1267;
        11'h4F4: data = 8'd1268;
        11'h4F5: data = 8'd1269;
        11'h4F6: data = 8'd1270;
        11'h4F7: data = 8'd1271;
        11'h4F8: data = 8'd1272;
        11'h4F9: data = 8'd1273;
        11'h4FA: data = 8'd1274;
        11'h4FB: data = 8'd1275;
        11'h4FC: data = 8'd1276;
        11'h4FD: data = 8'd1277;
        11'h4FE: data = 8'd1278;
        11'h4FF: data = 8'd1279;
        11'h500: data = 8'd1280;
        11'h501: data = 8'd1281;
        11'h502: data = 8'd1282;
        11'h503: data = 8'd1283;
        11'h504: data = 8'd1284;
        11'h505: data = 8'd1285;
        11'h506: data = 8'd1286;
        11'h507: data = 8'd1287;
        11'h508: data = 8'd1288;
        11'h509: data = 8'd1289;
        11'h50A: data = 8'd1290;
        11'h50B: data = 8'd1291;
        11'h50C: data = 8'd1292;
        11'h50D: data = 8'd1293;
        11'h50E: data = 8'd1294;
        11'h50F: data = 8'd1295;
        11'h510: data = 8'd1296;
        11'h511: data = 8'd1297;
        11'h512: data = 8'd1298;
        11'h513: data = 8'd1299;
        11'h514: data = 8'd1300;
        11'h515: data = 8'd1301;
        11'h516: data = 8'd1302;
        11'h517: data = 8'd1303;
        11'h518: data = 8'd1304;
        11'h519: data = 8'd1305;
        11'h51A: data = 8'd1306;
        11'h51B: data = 8'd1307;
        11'h51C: data = 8'd1308;
        11'h51D: data = 8'd1309;
        11'h51E: data = 8'd1310;
        11'h51F: data = 8'd1311;
        11'h520: data = 8'd1312;
        11'h521: data = 8'd1313;
        11'h522: data = 8'd1314;
        11'h523: data = 8'd1315;
        11'h524: data = 8'd1316;
        11'h525: data = 8'd1317;
        11'h526: data = 8'd1318;
        11'h527: data = 8'd1319;
        11'h528: data = 8'd1320;
        11'h529: data = 8'd1321;
        11'h52A: data = 8'd1322;
        11'h52B: data = 8'd1323;
        11'h52C: data = 8'd1324;
        11'h52D: data = 8'd1325;
        11'h52E: data = 8'd1326;
        11'h52F: data = 8'd1327;
        11'h530: data = 8'd1328;
        11'h531: data = 8'd1329;
        11'h532: data = 8'd1330;
        11'h533: data = 8'd1331;
        11'h534: data = 8'd1332;
        11'h535: data = 8'd1333;
        11'h536: data = 8'd1334;
        11'h537: data = 8'd1335;
        11'h538: data = 8'd1336;
        11'h539: data = 8'd1337;
        11'h53A: data = 8'd1338;
        11'h53B: data = 8'd1339;
        11'h53C: data = 8'd1340;
        11'h53D: data = 8'd1341;
        11'h53E: data = 8'd1342;
        11'h53F: data = 8'd1343;
        11'h540: data = 8'd1344;
        11'h541: data = 8'd1345;
        11'h542: data = 8'd1346;
        11'h543: data = 8'd1347;
        11'h544: data = 8'd1348;
        11'h545: data = 8'd1349;
        11'h546: data = 8'd1350;
        11'h547: data = 8'd1351;
        11'h548: data = 8'd1352;
        11'h549: data = 8'd1353;
        11'h54A: data = 8'd1354;
        11'h54B: data = 8'd1355;
        11'h54C: data = 8'd1356;
        11'h54D: data = 8'd1357;
        11'h54E: data = 8'd1358;
        11'h54F: data = 8'd1359;
        11'h550: data = 8'd1360;
        11'h551: data = 8'd1361;
        11'h552: data = 8'd1362;
        11'h553: data = 8'd1363;
        11'h554: data = 8'd1364;
        11'h555: data = 8'd1365;
        11'h556: data = 8'd1366;
        11'h557: data = 8'd1367;
        11'h558: data = 8'd1368;
        11'h559: data = 8'd1369;
        11'h55A: data = 8'd1370;
        11'h55B: data = 8'd1371;
        11'h55C: data = 8'd1372;
        11'h55D: data = 8'd1373;
        11'h55E: data = 8'd1374;
        11'h55F: data = 8'd1375;
        11'h560: data = 8'd1376;
        11'h561: data = 8'd1377;
        11'h562: data = 8'd1378;
        11'h563: data = 8'd1379;
        11'h564: data = 8'd1380;
        11'h565: data = 8'd1381;
        11'h566: data = 8'd1382;
        11'h567: data = 8'd1383;
        11'h568: data = 8'd1384;
        11'h569: data = 8'd1385;
        11'h56A: data = 8'd1386;
        11'h56B: data = 8'd1387;
        11'h56C: data = 8'd1388;
        11'h56D: data = 8'd1389;
        11'h56E: data = 8'd1390;
        11'h56F: data = 8'd1391;
        11'h570: data = 8'd1392;
        11'h571: data = 8'd1393;
        11'h572: data = 8'd1394;
        11'h573: data = 8'd1395;
        11'h574: data = 8'd1396;
        11'h575: data = 8'd1397;
        11'h576: data = 8'd1398;
        11'h577: data = 8'd1399;
        11'h578: data = 8'd1400;
        11'h579: data = 8'd1401;
        11'h57A: data = 8'd1402;
        11'h57B: data = 8'd1403;
        11'h57C: data = 8'd1404;
        11'h57D: data = 8'd1405;
        11'h57E: data = 8'd1406;
        11'h57F: data = 8'd1407;
        11'h580: data = 8'd1408;
        11'h581: data = 8'd1409;
        11'h582: data = 8'd1410;
        11'h583: data = 8'd1411;
        11'h584: data = 8'd1412;
        11'h585: data = 8'd1413;
        11'h586: data = 8'd1414;
        11'h587: data = 8'd1415;
        11'h588: data = 8'd1416;
        11'h589: data = 8'd1417;
        11'h58A: data = 8'd1418;
        11'h58B: data = 8'd1419;
        11'h58C: data = 8'd1420;
        11'h58D: data = 8'd1421;
        11'h58E: data = 8'd1422;
        11'h58F: data = 8'd1423;
        11'h590: data = 8'd1424;
        11'h591: data = 8'd1425;
        11'h592: data = 8'd1426;
        11'h593: data = 8'd1427;
        11'h594: data = 8'd1428;
        11'h595: data = 8'd1429;
        11'h596: data = 8'd1430;
        11'h597: data = 8'd1431;
        11'h598: data = 8'd1432;
        11'h599: data = 8'd1433;
        11'h59A: data = 8'd1434;
        11'h59B: data = 8'd1435;
        11'h59C: data = 8'd1436;
        11'h59D: data = 8'd1437;
        11'h59E: data = 8'd1438;
        11'h59F: data = 8'd1439;
        11'h5A0: data = 8'd1440;
        11'h5A1: data = 8'd1441;
        11'h5A2: data = 8'd1442;
        11'h5A3: data = 8'd1443;
        11'h5A4: data = 8'd1444;
        11'h5A5: data = 8'd1445;
        11'h5A6: data = 8'd1446;
        11'h5A7: data = 8'd1447;
        11'h5A8: data = 8'd1448;
        11'h5A9: data = 8'd1449;
        11'h5AA: data = 8'd1450;
        11'h5AB: data = 8'd1451;
        11'h5AC: data = 8'd1452;
        11'h5AD: data = 8'd1453;
        11'h5AE: data = 8'd1454;
        11'h5AF: data = 8'd1455;
        11'h5B0: data = 8'd1456;
        11'h5B1: data = 8'd1457;
        11'h5B2: data = 8'd1458;
        11'h5B3: data = 8'd1459;
        11'h5B4: data = 8'd1460;
        11'h5B5: data = 8'd1461;
        11'h5B6: data = 8'd1462;
        11'h5B7: data = 8'd1463;
        11'h5B8: data = 8'd1464;
        11'h5B9: data = 8'd1465;
        11'h5BA: data = 8'd1466;
        11'h5BB: data = 8'd1467;
        11'h5BC: data = 8'd1468;
        11'h5BD: data = 8'd1469;
        11'h5BE: data = 8'd1470;
        11'h5BF: data = 8'd1471;
        11'h5C0: data = 8'd1472;
        11'h5C1: data = 8'd1473;
        11'h5C2: data = 8'd1474;
        11'h5C3: data = 8'd1475;
        11'h5C4: data = 8'd1476;
        11'h5C5: data = 8'd1477;
        11'h5C6: data = 8'd1478;
        11'h5C7: data = 8'd1479;
        11'h5C8: data = 8'd1480;
        11'h5C9: data = 8'd1481;
        11'h5CA: data = 8'd1482;
        11'h5CB: data = 8'd1483;
        11'h5CC: data = 8'd1484;
        11'h5CD: data = 8'd1485;
        11'h5CE: data = 8'd1486;
        11'h5CF: data = 8'd1487;
        11'h5D0: data = 8'd1488;
        11'h5D1: data = 8'd1489;
        11'h5D2: data = 8'd1490;
        11'h5D3: data = 8'd1491;
        11'h5D4: data = 8'd1492;
        11'h5D5: data = 8'd1493;
        11'h5D6: data = 8'd1494;
        11'h5D7: data = 8'd1495;
        11'h5D8: data = 8'd1496;
        11'h5D9: data = 8'd1497;
        11'h5DA: data = 8'd1498;
        11'h5DB: data = 8'd1499;
        11'h5DC: data = 8'd1500;
        11'h5DD: data = 8'd1501;
        11'h5DE: data = 8'd1502;
        11'h5DF: data = 8'd1503;
        11'h5E0: data = 8'd1504;
        11'h5E1: data = 8'd1505;
        11'h5E2: data = 8'd1506;
        11'h5E3: data = 8'd1507;
        11'h5E4: data = 8'd1508;
        11'h5E5: data = 8'd1509;
        11'h5E6: data = 8'd1510;
        11'h5E7: data = 8'd1511;
        11'h5E8: data = 8'd1512;
        11'h5E9: data = 8'd1513;
        11'h5EA: data = 8'd1514;
        11'h5EB: data = 8'd1515;
        11'h5EC: data = 8'd1516;
        11'h5ED: data = 8'd1517;
        11'h5EE: data = 8'd1518;
        11'h5EF: data = 8'd1519;
        11'h5F0: data = 8'd1520;
        11'h5F1: data = 8'd1521;
        11'h5F2: data = 8'd1522;
        11'h5F3: data = 8'd1523;
        11'h5F4: data = 8'd1524;
        11'h5F5: data = 8'd1525;
        11'h5F6: data = 8'd1526;
        11'h5F7: data = 8'd1527;
        11'h5F8: data = 8'd1528;
        11'h5F9: data = 8'd1529;
        11'h5FA: data = 8'd1530;
        11'h5FB: data = 8'd1531;
        11'h5FC: data = 8'd1532;
        11'h5FD: data = 8'd1533;
        11'h5FE: data = 8'd1534;
        11'h5FF: data = 8'd1535;
        11'h600: data = 8'd1536;
        11'h601: data = 8'd1537;
        11'h602: data = 8'd1538;
        11'h603: data = 8'd1539;
        11'h604: data = 8'd1540;
        11'h605: data = 8'd1541;
        11'h606: data = 8'd1542;
        11'h607: data = 8'd1543;
        11'h608: data = 8'd1544;
        11'h609: data = 8'd1545;
        11'h60A: data = 8'd1546;
        11'h60B: data = 8'd1547;
        11'h60C: data = 8'd1548;
        11'h60D: data = 8'd1549;
        11'h60E: data = 8'd1550;
        11'h60F: data = 8'd1551;
        11'h610: data = 8'd1552;
        11'h611: data = 8'd1553;
        11'h612: data = 8'd1554;
        11'h613: data = 8'd1555;
        11'h614: data = 8'd1556;
        11'h615: data = 8'd1557;
        11'h616: data = 8'd1558;
        11'h617: data = 8'd1559;
        11'h618: data = 8'd1560;
        11'h619: data = 8'd1561;
        11'h61A: data = 8'd1562;
        11'h61B: data = 8'd1563;
        11'h61C: data = 8'd1564;
        11'h61D: data = 8'd1565;
        11'h61E: data = 8'd1566;
        11'h61F: data = 8'd1567;
        11'h620: data = 8'd1568;
        11'h621: data = 8'd1569;
        11'h622: data = 8'd1570;
        11'h623: data = 8'd1571;
        11'h624: data = 8'd1572;
        11'h625: data = 8'd1573;
        11'h626: data = 8'd1574;
        11'h627: data = 8'd1575;
        11'h628: data = 8'd1576;
        11'h629: data = 8'd1577;
        11'h62A: data = 8'd1578;
        11'h62B: data = 8'd1579;
        11'h62C: data = 8'd1580;
        11'h62D: data = 8'd1581;
        11'h62E: data = 8'd1582;
        11'h62F: data = 8'd1583;
        11'h630: data = 8'd1584;
        11'h631: data = 8'd1585;
        11'h632: data = 8'd1586;
        11'h633: data = 8'd1587;
        11'h634: data = 8'd1588;
        11'h635: data = 8'd1589;
        11'h636: data = 8'd1590;
        11'h637: data = 8'd1591;
        11'h638: data = 8'd1592;
        11'h639: data = 8'd1593;
        11'h63A: data = 8'd1594;
        11'h63B: data = 8'd1595;
        11'h63C: data = 8'd1596;
        11'h63D: data = 8'd1597;
        11'h63E: data = 8'd1598;
        11'h63F: data = 8'd1599;
        11'h640: data = 8'd1600;
        11'h641: data = 8'd1601;
        11'h642: data = 8'd1602;
        11'h643: data = 8'd1603;
        11'h644: data = 8'd1604;
        11'h645: data = 8'd1605;
        11'h646: data = 8'd1606;
        11'h647: data = 8'd1607;
        11'h648: data = 8'd1608;
        11'h649: data = 8'd1609;
        11'h64A: data = 8'd1610;
        11'h64B: data = 8'd1611;
        11'h64C: data = 8'd1612;
        11'h64D: data = 8'd1613;
        11'h64E: data = 8'd1614;
        11'h64F: data = 8'd1615;
        11'h650: data = 8'd1616;
        11'h651: data = 8'd1617;
        11'h652: data = 8'd1618;
        11'h653: data = 8'd1619;
        11'h654: data = 8'd1620;
        11'h655: data = 8'd1621;
        11'h656: data = 8'd1622;
        11'h657: data = 8'd1623;
        11'h658: data = 8'd1624;
        11'h659: data = 8'd1625;
        11'h65A: data = 8'd1626;
        11'h65B: data = 8'd1627;
        11'h65C: data = 8'd1628;
        11'h65D: data = 8'd1629;
        11'h65E: data = 8'd1630;
        11'h65F: data = 8'd1631;
        11'h660: data = 8'd1632;
        11'h661: data = 8'd1633;
        11'h662: data = 8'd1634;
        11'h663: data = 8'd1635;
        11'h664: data = 8'd1636;
        11'h665: data = 8'd1637;
        11'h666: data = 8'd1638;
        11'h667: data = 8'd1639;
        11'h668: data = 8'd1640;
        11'h669: data = 8'd1641;
        11'h66A: data = 8'd1642;
        11'h66B: data = 8'd1643;
        11'h66C: data = 8'd1644;
        11'h66D: data = 8'd1645;
        11'h66E: data = 8'd1646;
        11'h66F: data = 8'd1647;
        11'h670: data = 8'd1648;
        11'h671: data = 8'd1649;
        11'h672: data = 8'd1650;
        11'h673: data = 8'd1651;
        11'h674: data = 8'd1652;
        11'h675: data = 8'd1653;
        11'h676: data = 8'd1654;
        11'h677: data = 8'd1655;
        11'h678: data = 8'd1656;
        11'h679: data = 8'd1657;
        11'h67A: data = 8'd1658;
        11'h67B: data = 8'd1659;
        11'h67C: data = 8'd1660;
        11'h67D: data = 8'd1661;
        11'h67E: data = 8'd1662;
        11'h67F: data = 8'd1663;
        11'h680: data = 8'd1664;
        11'h681: data = 8'd1665;
        11'h682: data = 8'd1666;
        11'h683: data = 8'd1667;
        11'h684: data = 8'd1668;
        11'h685: data = 8'd1669;
        11'h686: data = 8'd1670;
        11'h687: data = 8'd1671;
        11'h688: data = 8'd1672;
        11'h689: data = 8'd1673;
        11'h68A: data = 8'd1674;
        11'h68B: data = 8'd1675;
        11'h68C: data = 8'd1676;
        11'h68D: data = 8'd1677;
        11'h68E: data = 8'd1678;
        11'h68F: data = 8'd1679;
        11'h690: data = 8'd1680;
        11'h691: data = 8'd1681;
        11'h692: data = 8'd1682;
        11'h693: data = 8'd1683;
        11'h694: data = 8'd1684;
        11'h695: data = 8'd1685;
        11'h696: data = 8'd1686;
        11'h697: data = 8'd1687;
        11'h698: data = 8'd1688;
        11'h699: data = 8'd1689;
        11'h69A: data = 8'd1690;
        11'h69B: data = 8'd1691;
        11'h69C: data = 8'd1692;
        11'h69D: data = 8'd1693;
        11'h69E: data = 8'd1694;
        11'h69F: data = 8'd1695;
        11'h6A0: data = 8'd1696;
        11'h6A1: data = 8'd1697;
        11'h6A2: data = 8'd1698;
        11'h6A3: data = 8'd1699;
        11'h6A4: data = 8'd1700;
        11'h6A5: data = 8'd1701;
        11'h6A6: data = 8'd1702;
        11'h6A7: data = 8'd1703;
        11'h6A8: data = 8'd1704;
        11'h6A9: data = 8'd1705;
        11'h6AA: data = 8'd1706;
        11'h6AB: data = 8'd1707;
        11'h6AC: data = 8'd1708;
        11'h6AD: data = 8'd1709;
        11'h6AE: data = 8'd1710;
        11'h6AF: data = 8'd1711;
        11'h6B0: data = 8'd1712;
        11'h6B1: data = 8'd1713;
        11'h6B2: data = 8'd1714;
        11'h6B3: data = 8'd1715;
        11'h6B4: data = 8'd1716;
        11'h6B5: data = 8'd1717;
        11'h6B6: data = 8'd1718;
        11'h6B7: data = 8'd1719;
        11'h6B8: data = 8'd1720;
        11'h6B9: data = 8'd1721;
        11'h6BA: data = 8'd1722;
        11'h6BB: data = 8'd1723;
        11'h6BC: data = 8'd1724;
        11'h6BD: data = 8'd1725;
        11'h6BE: data = 8'd1726;
        11'h6BF: data = 8'd1727;
        11'h6C0: data = 8'd1728;
        11'h6C1: data = 8'd1729;
        11'h6C2: data = 8'd1730;
        11'h6C3: data = 8'd1731;
        11'h6C4: data = 8'd1732;
        11'h6C5: data = 8'd1733;
        11'h6C6: data = 8'd1734;
        11'h6C7: data = 8'd1735;
        11'h6C8: data = 8'd1736;
        11'h6C9: data = 8'd1737;
        11'h6CA: data = 8'd1738;
        11'h6CB: data = 8'd1739;
        11'h6CC: data = 8'd1740;
        11'h6CD: data = 8'd1741;
        11'h6CE: data = 8'd1742;
        11'h6CF: data = 8'd1743;
        11'h6D0: data = 8'd1744;
        11'h6D1: data = 8'd1745;
        11'h6D2: data = 8'd1746;
        11'h6D3: data = 8'd1747;
        11'h6D4: data = 8'd1748;
        11'h6D5: data = 8'd1749;
        11'h6D6: data = 8'd1750;
        11'h6D7: data = 8'd1751;
        11'h6D8: data = 8'd1752;
        11'h6D9: data = 8'd1753;
        11'h6DA: data = 8'd1754;
        11'h6DB: data = 8'd1755;
        11'h6DC: data = 8'd1756;
        11'h6DD: data = 8'd1757;
        11'h6DE: data = 8'd1758;
        11'h6DF: data = 8'd1759;
        11'h6E0: data = 8'd1760;
        11'h6E1: data = 8'd1761;
        11'h6E2: data = 8'd1762;
        11'h6E3: data = 8'd1763;
        11'h6E4: data = 8'd1764;
        11'h6E5: data = 8'd1765;
        11'h6E6: data = 8'd1766;
        11'h6E7: data = 8'd1767;
        11'h6E8: data = 8'd1768;
        11'h6E9: data = 8'd1769;
        11'h6EA: data = 8'd1770;
        11'h6EB: data = 8'd1771;
        11'h6EC: data = 8'd1772;
        11'h6ED: data = 8'd1773;
        11'h6EE: data = 8'd1774;
        11'h6EF: data = 8'd1775;
        11'h6F0: data = 8'd1776;
        11'h6F1: data = 8'd1777;
        11'h6F2: data = 8'd1778;
        11'h6F3: data = 8'd1779;
        11'h6F4: data = 8'd1780;
        11'h6F5: data = 8'd1781;
        11'h6F6: data = 8'd1782;
        11'h6F7: data = 8'd1783;
        11'h6F8: data = 8'd1784;
        11'h6F9: data = 8'd1785;
        11'h6FA: data = 8'd1786;
        11'h6FB: data = 8'd1787;
        11'h6FC: data = 8'd1788;
        11'h6FD: data = 8'd1789;
        11'h6FE: data = 8'd1790;
        11'h6FF: data = 8'd1791;
        11'h700: data = 8'd1792;
        11'h701: data = 8'd1793;
        11'h702: data = 8'd1794;
        11'h703: data = 8'd1795;
        11'h704: data = 8'd1796;
        11'h705: data = 8'd1797;
        11'h706: data = 8'd1798;
        11'h707: data = 8'd1799;
        11'h708: data = 8'd1800;
        11'h709: data = 8'd1801;
        11'h70A: data = 8'd1802;
        11'h70B: data = 8'd1803;
        11'h70C: data = 8'd1804;
        11'h70D: data = 8'd1805;
        11'h70E: data = 8'd1806;
        11'h70F: data = 8'd1807;
        11'h710: data = 8'd1808;
        11'h711: data = 8'd1809;
        11'h712: data = 8'd1810;
        11'h713: data = 8'd1811;
        11'h714: data = 8'd1812;
        11'h715: data = 8'd1813;
        11'h716: data = 8'd1814;
        11'h717: data = 8'd1815;
        11'h718: data = 8'd1816;
        11'h719: data = 8'd1817;
        11'h71A: data = 8'd1818;
        11'h71B: data = 8'd1819;
        11'h71C: data = 8'd1820;
        11'h71D: data = 8'd1821;
        11'h71E: data = 8'd1822;
        11'h71F: data = 8'd1823;
        11'h720: data = 8'd1824;
        11'h721: data = 8'd1825;
        11'h722: data = 8'd1826;
        11'h723: data = 8'd1827;
        11'h724: data = 8'd1828;
        11'h725: data = 8'd1829;
        11'h726: data = 8'd1830;
        11'h727: data = 8'd1831;
        11'h728: data = 8'd1832;
        11'h729: data = 8'd1833;
        11'h72A: data = 8'd1834;
        11'h72B: data = 8'd1835;
        11'h72C: data = 8'd1836;
        11'h72D: data = 8'd1837;
        11'h72E: data = 8'd1838;
        11'h72F: data = 8'd1839;
        11'h730: data = 8'd1840;
        11'h731: data = 8'd1841;
        11'h732: data = 8'd1842;
        11'h733: data = 8'd1843;
        11'h734: data = 8'd1844;
        11'h735: data = 8'd1845;
        11'h736: data = 8'd1846;
        11'h737: data = 8'd1847;
        11'h738: data = 8'd1848;
        11'h739: data = 8'd1849;
        11'h73A: data = 8'd1850;
        11'h73B: data = 8'd1851;
        11'h73C: data = 8'd1852;
        11'h73D: data = 8'd1853;
        11'h73E: data = 8'd1854;
        11'h73F: data = 8'd1855;
        11'h740: data = 8'd1856;
        11'h741: data = 8'd1857;
        11'h742: data = 8'd1858;
        11'h743: data = 8'd1859;
        11'h744: data = 8'd1860;
        11'h745: data = 8'd1861;
        11'h746: data = 8'd1862;
        11'h747: data = 8'd1863;
        11'h748: data = 8'd1864;
        11'h749: data = 8'd1865;
        11'h74A: data = 8'd1866;
        11'h74B: data = 8'd1867;
        11'h74C: data = 8'd1868;
        11'h74D: data = 8'd1869;
        11'h74E: data = 8'd1870;
        11'h74F: data = 8'd1871;
        11'h750: data = 8'd1872;
        11'h751: data = 8'd1873;
        11'h752: data = 8'd1874;
        11'h753: data = 8'd1875;
        11'h754: data = 8'd1876;
        11'h755: data = 8'd1877;
        11'h756: data = 8'd1878;
        11'h757: data = 8'd1879;
        11'h758: data = 8'd1880;
        11'h759: data = 8'd1881;
        11'h75A: data = 8'd1882;
        11'h75B: data = 8'd1883;
        11'h75C: data = 8'd1884;
        11'h75D: data = 8'd1885;
        11'h75E: data = 8'd1886;
        11'h75F: data = 8'd1887;
        11'h760: data = 8'd1888;
        11'h761: data = 8'd1889;
        11'h762: data = 8'd1890;
        11'h763: data = 8'd1891;
        11'h764: data = 8'd1892;
        11'h765: data = 8'd1893;
        11'h766: data = 8'd1894;
        11'h767: data = 8'd1895;
        11'h768: data = 8'd1896;
        11'h769: data = 8'd1897;
        11'h76A: data = 8'd1898;
        11'h76B: data = 8'd1899;
        11'h76C: data = 8'd1900;
        11'h76D: data = 8'd1901;
        11'h76E: data = 8'd1902;
        11'h76F: data = 8'd1903;
        11'h770: data = 8'd1904;
        11'h771: data = 8'd1905;
        11'h772: data = 8'd1906;
        11'h773: data = 8'd1907;
        11'h774: data = 8'd1908;
        11'h775: data = 8'd1909;
        11'h776: data = 8'd1910;
        11'h777: data = 8'd1911;
        11'h778: data = 8'd1912;
        11'h779: data = 8'd1913;
        11'h77A: data = 8'd1914;
        11'h77B: data = 8'd1915;
        11'h77C: data = 8'd1916;
        11'h77D: data = 8'd1917;
        11'h77E: data = 8'd1918;
        11'h77F: data = 8'd1919;
        11'h780: data = 8'd1920;
        11'h781: data = 8'd1921;
        11'h782: data = 8'd1922;
        11'h783: data = 8'd1923;
        11'h784: data = 8'd1924;
        11'h785: data = 8'd1925;
        11'h786: data = 8'd1926;
        11'h787: data = 8'd1927;
        11'h788: data = 8'd1928;
        11'h789: data = 8'd1929;
        11'h78A: data = 8'd1930;
        11'h78B: data = 8'd1931;
        11'h78C: data = 8'd1932;
        11'h78D: data = 8'd1933;
        11'h78E: data = 8'd1934;
        11'h78F: data = 8'd1935;
        11'h790: data = 8'd1936;
        11'h791: data = 8'd1937;
        11'h792: data = 8'd1938;
        11'h793: data = 8'd1939;
        11'h794: data = 8'd1940;
        11'h795: data = 8'd1941;
        11'h796: data = 8'd1942;
        11'h797: data = 8'd1943;
        11'h798: data = 8'd1944;
        11'h799: data = 8'd1945;
        11'h79A: data = 8'd1946;
        11'h79B: data = 8'd1947;
        11'h79C: data = 8'd1948;
        11'h79D: data = 8'd1949;
        11'h79E: data = 8'd1950;
        11'h79F: data = 8'd1951;
        11'h7A0: data = 8'd1952;
        11'h7A1: data = 8'd1953;
        11'h7A2: data = 8'd1954;
        11'h7A3: data = 8'd1955;
        11'h7A4: data = 8'd1956;
        11'h7A5: data = 8'd1957;
        11'h7A6: data = 8'd1958;
        11'h7A7: data = 8'd1959;
        11'h7A8: data = 8'd1960;
        11'h7A9: data = 8'd1961;
        11'h7AA: data = 8'd1962;
        11'h7AB: data = 8'd1963;
        11'h7AC: data = 8'd1964;
        11'h7AD: data = 8'd1965;
        11'h7AE: data = 8'd1966;
        11'h7AF: data = 8'd1967;
        11'h7B0: data = 8'd1968;
        11'h7B1: data = 8'd1969;
        11'h7B2: data = 8'd1970;
        11'h7B3: data = 8'd1971;
        11'h7B4: data = 8'd1972;
        11'h7B5: data = 8'd1973;
        11'h7B6: data = 8'd1974;
        11'h7B7: data = 8'd1975;
        11'h7B8: data = 8'd1976;
        11'h7B9: data = 8'd1977;
        11'h7BA: data = 8'd1978;
        11'h7BB: data = 8'd1979;
        11'h7BC: data = 8'd1980;
        11'h7BD: data = 8'd1981;
        11'h7BE: data = 8'd1982;
        11'h7BF: data = 8'd1983;
        11'h7C0: data = 8'd1984;
        11'h7C1: data = 8'd1985;
        11'h7C2: data = 8'd1986;
        11'h7C3: data = 8'd1987;
        11'h7C4: data = 8'd1988;
        11'h7C5: data = 8'd1989;
        11'h7C6: data = 8'd1990;
        11'h7C7: data = 8'd1991;
        11'h7C8: data = 8'd1992;
        11'h7C9: data = 8'd1993;
        11'h7CA: data = 8'd1994;
        11'h7CB: data = 8'd1995;
        11'h7CC: data = 8'd1996;
        11'h7CD: data = 8'd1997;
        11'h7CE: data = 8'd1998;
        11'h7CF: data = 8'd1999;
        11'h7D0: data = 8'd2000;
        11'h7D1: data = 8'd2001;
        11'h7D2: data = 8'd2002;
        11'h7D3: data = 8'd2003;
        11'h7D4: data = 8'd2004;
        11'h7D5: data = 8'd2005;
        11'h7D6: data = 8'd2006;
        11'h7D7: data = 8'd2007;
        11'h7D8: data = 8'd2008;
        11'h7D9: data = 8'd2009;
        11'h7DA: data = 8'd2010;
        11'h7DB: data = 8'd2011;
        11'h7DC: data = 8'd2012;
        11'h7DD: data = 8'd2013;
        11'h7DE: data = 8'd2014;
        11'h7DF: data = 8'd2015;
        11'h7E0: data = 8'd2016;
        11'h7E1: data = 8'd2017;
        11'h7E2: data = 8'd2018;
        11'h7E3: data = 8'd2019;
        11'h7E4: data = 8'd2020;
        11'h7E5: data = 8'd2021;
        11'h7E6: data = 8'd2022;
        11'h7E7: data = 8'd2023;
        11'h7E8: data = 8'd2024;
        11'h7E9: data = 8'd2025;
        11'h7EA: data = 8'd2026;
        11'h7EB: data = 8'd2027;
        11'h7EC: data = 8'd2028;
        11'h7ED: data = 8'd2029;
        11'h7EE: data = 8'd2030;
        11'h7EF: data = 8'd2031;
        11'h7F0: data = 8'd2032;
        11'h7F1: data = 8'd2033;
        11'h7F2: data = 8'd2034;
        11'h7F3: data = 8'd2035;
        11'h7F4: data = 8'd2036;
        11'h7F5: data = 8'd2037;
        11'h7F6: data = 8'd2038;
        11'h7F7: data = 8'd2039;
        11'h7F8: data = 8'd2040;
        11'h7F9: data = 8'd2041;
        11'h7FA: data = 8'd2042;
        11'h7FB: data = 8'd2043;
        11'h7FC: data = 8'd2044;
        11'h7FD: data = 8'd2045;
        11'h7FE: data = 8'd2046;
        11'h7FF: data = 8'd2047;
        default: data = '0;
    endcase
end


    

endmodule

